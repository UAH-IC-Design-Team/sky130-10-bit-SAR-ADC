magic
tech sky130A
timestamp 1668278360
<< metal4 >>
rect -17250 12750 -5200 12900
rect -17250 12500 -17200 12750
rect -16450 12500 -16400 12750
rect -15650 12500 -15600 12750
rect -14850 12500 -14800 12750
rect -14050 12500 -14000 12750
rect -13250 12500 -13200 12750
rect -12450 12500 -12400 12750
rect -11650 12500 -11600 12750
rect -10850 12500 -10800 12750
rect -10050 12500 -10000 12750
rect -9250 12500 -9200 12750
rect -8450 12500 -8400 12750
rect -7650 12500 -7600 12750
rect -6850 12500 -6800 12750
rect -6050 12500 -6000 12750
rect -5250 12500 -5200 12750
rect -4450 12750 1200 12900
rect -4450 12500 -4400 12750
rect -3650 12500 -3600 12750
rect -2850 12500 -2800 12750
rect -2050 12500 -2000 12750
rect -1250 12500 -1200 12750
rect -450 12500 -400 12750
rect 350 12500 400 12750
rect 1150 12500 1200 12750
rect 1950 12750 14000 12900
rect 1950 12500 2000 12750
rect 2750 12500 2800 12750
rect 3550 12500 3600 12750
rect 4350 12500 4400 12750
rect 5150 12500 5200 12750
rect 5950 12500 6000 12750
rect 6750 12500 6800 12750
rect 7550 12500 7600 12750
rect 8350 12500 8400 12750
rect 9150 12500 9200 12750
rect 9950 12500 10000 12750
rect 10750 12500 10800 12750
rect 11550 12500 11600 12750
rect 12350 12500 12400 12750
rect 13150 12500 13200 12750
rect 13950 12500 14000 12750
rect 14750 12750 20400 12900
rect 14750 12500 14800 12750
rect 15550 12500 15600 12750
rect 16350 12500 16400 12750
rect 17150 12500 17200 12750
rect 17950 12500 18000 12750
rect 18750 12500 18800 12750
rect 19550 12500 19600 12750
rect 20350 12500 20400 12750
rect 21150 12750 23600 12900
rect 21150 12500 21200 12750
rect 21950 12500 22000 12750
rect 22750 12500 22800 12750
rect 23550 12500 23600 12750
rect 24350 12750 25200 12900
rect 24350 12500 24400 12750
rect 25150 12500 25200 12750
rect 25950 12500 26000 12900
rect 26750 12750 29200 12900
rect 26750 12500 26800 12750
rect 27550 12500 27600 12750
rect 28350 12500 28400 12750
rect 29150 12500 29200 12750
rect 29950 12750 30800 12900
rect 29950 12500 30000 12750
rect 30750 12500 30800 12750
rect 31550 12500 31600 12900
rect 32350 7150 34800 7300
rect 32350 7100 32400 7150
rect 33150 7100 33200 7150
rect 33950 7100 34000 7150
rect 34750 7100 34800 7150
rect 35550 7150 36400 7300
rect 35550 7100 35600 7150
rect 36350 7100 36400 7150
rect 37150 7100 37200 7300
rect 37950 7150 40400 7300
rect 37950 7100 38000 7150
rect 38750 7100 38800 7150
rect 39550 7100 39600 7150
rect 40350 7100 40400 7150
rect 41150 7150 42000 7300
rect 41150 7100 41200 7150
rect 41950 7100 42000 7150
rect 42750 7100 42800 7300
rect 43550 7100 43600 7300
rect -16910 6450 -16850 6500
rect -16110 6450 -16050 6500
rect -15310 6450 -15250 6500
rect -14510 6450 -14450 6500
rect -13710 6450 -13650 6500
rect -12910 6450 -12850 6500
rect -12110 6450 -12050 6500
rect -11310 6450 -11250 6500
rect -10510 6450 -10450 6500
rect -9710 6450 -9650 6500
rect -8910 6450 -8850 6500
rect -8110 6450 -8050 6500
rect -7310 6450 -7250 6500
rect -6510 6450 -6450 6500
rect -5710 6450 -5650 6500
rect -4910 6450 -4850 6500
rect -4110 6450 -4050 6500
rect -3310 6450 -3250 6500
rect -2510 6450 -2450 6500
rect -1710 6450 -1650 6500
rect -910 6450 -850 6500
rect -110 6450 -50 6500
rect 690 6450 750 6500
rect 1490 6450 1550 6500
rect 2290 6450 2350 6500
rect 3090 6450 3150 6500
rect 3890 6450 3950 6500
rect 4690 6450 4750 6500
rect 5490 6450 5550 6500
rect 6290 6450 6350 6500
rect 7090 6450 7150 6500
rect 7890 6450 7950 6500
rect 8690 6450 8750 6500
rect 9490 6450 9550 6500
rect 10290 6450 10350 6500
rect 11090 6450 11150 6500
rect 11890 6450 11950 6500
rect 12690 6450 12750 6500
rect 13490 6450 13550 6500
rect 14290 6450 14350 6500
rect 15090 6450 15150 6500
rect 15890 6450 15950 6500
rect 16690 6450 16750 6500
rect 17490 6450 17550 6500
rect 18290 6450 18350 6500
rect 19090 6450 19150 6500
rect 19890 6450 19950 6500
rect 20690 6450 20750 6500
rect 21490 6450 21550 6500
rect 22290 6450 22350 6500
rect 23090 6450 23150 6500
rect 23890 6450 23950 6500
rect 24690 6450 24750 6500
rect 25490 6450 25550 6500
rect 26290 6450 26350 6500
rect 27090 6450 27150 6500
rect 27890 6450 27950 6500
rect 28690 6450 28750 6500
rect 29490 6450 29550 6500
rect 30290 6450 30350 6500
rect 31090 6450 31150 6500
rect 31890 6450 31950 6500
rect 32690 6450 32750 6500
rect 33490 6450 33550 6500
rect 34290 6450 34350 6500
rect 35090 6450 35150 6500
rect 35890 6450 35950 6500
rect 36690 6450 36750 6500
rect 37490 6450 37550 6500
rect 38290 6450 38350 6500
rect 39090 6450 39150 6500
rect 39890 6450 39950 6500
rect 40690 6450 40750 6500
rect 41490 6450 41550 6500
rect 42290 6450 42350 6500
rect 43090 6450 43150 6500
rect 43890 6450 43950 6500
rect -16910 6250 43950 6450
rect -16910 4950 43950 5150
rect -16910 4900 -16850 4950
rect -16110 4900 -16050 4950
rect -15310 4900 -15250 4950
rect -14510 4900 -14450 4950
rect -13710 4900 -13650 4950
rect -12910 4900 -12850 4950
rect -12110 4900 -12050 4950
rect -11310 4900 -11250 4950
rect -10510 4900 -10450 4950
rect -9710 4900 -9650 4950
rect -8910 4900 -8850 4950
rect -8110 4900 -8050 4950
rect -7310 4900 -7250 4950
rect -6510 4900 -6450 4950
rect -5710 4900 -5650 4950
rect -4910 4900 -4850 4950
rect -4110 4900 -4050 4950
rect -3310 4900 -3250 4950
rect -2510 4900 -2450 4950
rect -1710 4900 -1650 4950
rect -910 4900 -850 4950
rect -110 4900 -50 4950
rect 690 4900 750 4950
rect 1490 4900 1550 4950
rect 2290 4900 2350 4950
rect 3090 4900 3150 4950
rect 3890 4900 3950 4950
rect 4690 4900 4750 4950
rect 5490 4900 5550 4950
rect 6290 4900 6350 4950
rect 7090 4900 7150 4950
rect 7890 4900 7950 4950
rect 8690 4900 8750 4950
rect 9490 4900 9550 4950
rect 10290 4900 10350 4950
rect 11090 4900 11150 4950
rect 11890 4900 11950 4950
rect 12690 4900 12750 4950
rect 13490 4900 13550 4950
rect 14290 4900 14350 4950
rect 15090 4900 15150 4950
rect 15890 4900 15950 4950
rect 16690 4900 16750 4950
rect 17490 4900 17550 4950
rect 18290 4900 18350 4950
rect 19090 4900 19150 4950
rect 19890 4900 19950 4950
rect 20690 4900 20750 4950
rect 21490 4900 21550 4950
rect 22290 4900 22350 4950
rect 23090 4900 23150 4950
rect 23890 4900 23950 4950
rect 24690 4900 24750 4950
rect 25490 4900 25550 4950
rect 26290 4900 26350 4950
rect 27090 4900 27150 4950
rect 27890 4900 27950 4950
rect 28690 4900 28750 4950
rect 29490 4900 29550 4950
rect 30290 4900 30350 4950
rect 31090 4900 31150 4950
rect 31890 4900 31950 4950
rect 32690 4900 32750 4950
rect 33490 4900 33550 4950
rect 34290 4900 34350 4950
rect 35090 4900 35150 4950
rect 35890 4900 35950 4950
rect 36690 4900 36750 4950
rect 37490 4900 37550 4950
rect 38290 4900 38350 4950
rect 39090 4900 39150 4950
rect 39890 4900 39950 4950
rect 40690 4900 40750 4950
rect 41490 4900 41550 4950
rect 42290 4900 42350 4950
rect 43090 4900 43150 4950
rect 43890 4900 43950 4950
rect 32350 4250 32400 4300
rect 33150 4250 33200 4300
rect 33950 4250 34000 4300
rect 34750 4250 34800 4300
rect 32350 4100 34800 4250
rect 35550 4250 35600 4300
rect 36350 4250 36400 4300
rect 35550 4100 36400 4250
rect 37150 4100 37200 4300
rect 37950 4250 38000 4300
rect 38750 4250 38800 4300
rect 39550 4250 39600 4300
rect 40350 4250 40400 4300
rect 37950 4100 40400 4250
rect 41150 4250 41200 4300
rect 41950 4250 42000 4300
rect 41150 4100 42000 4250
rect 42750 4100 42800 4300
rect 43550 4100 43600 4300
rect -17250 -1350 -17200 -1100
rect -16450 -1350 -16400 -1100
rect -15650 -1350 -15600 -1100
rect -14850 -1350 -14800 -1100
rect -14050 -1350 -14000 -1100
rect -13250 -1350 -13200 -1100
rect -12450 -1350 -12400 -1100
rect -11650 -1350 -11600 -1100
rect -10850 -1350 -10800 -1100
rect -10050 -1350 -10000 -1100
rect -9250 -1350 -9200 -1100
rect -8450 -1350 -8400 -1100
rect -7650 -1350 -7600 -1100
rect -6850 -1350 -6800 -1100
rect -6050 -1350 -6000 -1100
rect -5250 -1350 -5200 -1100
rect -17250 -1500 -5200 -1350
rect -4450 -1350 -4400 -1100
rect -3650 -1350 -3600 -1100
rect -2850 -1350 -2800 -1100
rect -2050 -1350 -2000 -1100
rect -1250 -1350 -1200 -1100
rect -450 -1350 -400 -1100
rect 350 -1350 400 -1100
rect 1150 -1350 1200 -1100
rect -4450 -1500 1200 -1350
rect 1950 -1350 2000 -1100
rect 2750 -1350 2800 -1100
rect 3550 -1350 3600 -1100
rect 4350 -1350 4400 -1100
rect 5150 -1350 5200 -1100
rect 5950 -1350 6000 -1100
rect 6750 -1350 6800 -1100
rect 7550 -1350 7600 -1100
rect 8350 -1350 8400 -1100
rect 9150 -1350 9200 -1100
rect 9950 -1350 10000 -1100
rect 10750 -1350 10800 -1100
rect 11550 -1350 11600 -1100
rect 12350 -1350 12400 -1100
rect 13150 -1350 13200 -1100
rect 13950 -1350 14000 -1100
rect 1950 -1500 14000 -1350
rect 14750 -1350 14800 -1100
rect 15550 -1350 15600 -1100
rect 16350 -1350 16400 -1100
rect 17150 -1350 17200 -1100
rect 17950 -1350 18000 -1100
rect 18750 -1350 18800 -1100
rect 19550 -1350 19600 -1100
rect 20350 -1350 20400 -1100
rect 14750 -1500 20400 -1350
rect 21150 -1350 21200 -1100
rect 21950 -1350 22000 -1100
rect 22750 -1350 22800 -1100
rect 23550 -1350 23600 -1100
rect 21150 -1500 23600 -1350
rect 24350 -1350 24400 -1100
rect 25150 -1350 25200 -1100
rect 24350 -1500 25200 -1350
rect 25950 -1500 26000 -1100
rect 26750 -1350 26800 -1100
rect 27550 -1350 27600 -1100
rect 28350 -1350 28400 -1100
rect 29150 -1350 29200 -1100
rect 26750 -1500 29200 -1350
rect 29950 -1350 30000 -1100
rect 30750 -1350 30800 -1100
rect 29950 -1500 30800 -1350
rect 31550 -1500 31600 -1100
use cap1  cap1_0
timestamp 1667663783
transform 1 0 36900 0 1 6500
box 0 0 650 600
use cap1  cap1_1
timestamp 1667663783
transform 1 0 42500 0 -1 4900
box 0 0 650 600
use cap1  cap1_2
timestamp 1667663783
transform 1 0 43300 0 -1 4900
box 0 0 650 600
use cap1  cap1_3
timestamp 1667663783
transform 1 0 36900 0 -1 4900
box 0 0 650 600
use cap1  cap1_4
timestamp 1667663783
transform 1 0 43300 0 1 6500
box 0 0 650 600
use cap1  cap1_5
timestamp 1667663783
transform 1 0 42500 0 1 6500
box 0 0 650 600
use cap2  cap2_0
timestamp 1667663783
transform 1 0 35300 0 1 6500
box 0 0 1450 600
use cap2  cap2_1
timestamp 1667663783
transform 1 0 40900 0 -1 4900
box 0 0 1450 600
use cap2  cap2_2
timestamp 1667663783
transform 1 0 35300 0 -1 4900
box 0 0 1450 600
use cap2  cap2_3
timestamp 1667663783
transform 1 0 40900 0 1 6500
box 0 0 1450 600
use cap4  cap4_0
timestamp 1667663783
transform 1 0 32100 0 1 6500
box 0 0 3050 600
use cap4  cap4_1
timestamp 1667663783
transform 1 0 37700 0 1 6500
box 0 0 3050 600
use cap4  cap4_2
timestamp 1667663783
transform 1 0 37700 0 -1 4900
box 0 0 3050 600
use cap4  cap4_3
timestamp 1667663783
transform 1 0 32100 0 -1 4900
box 0 0 3050 600
use cap8  cap8_0
timestamp 1667684479
transform 1 0 25700 0 1 6500
box 0 0 650 6200
use cap8  cap8_1
timestamp 1667684479
transform 1 0 31300 0 1 6500
box 0 0 650 6200
use cap8  cap8_2
timestamp 1667684479
transform 1 0 31300 0 -1 4900
box 0 0 650 6200
use cap8  cap8_3
timestamp 1667684479
transform 1 0 25700 0 -1 4900
box 0 0 650 6200
use cap16  cap16_0
timestamp 1667684462
transform 1 0 24100 0 1 6500
box 0 0 1450 6200
use cap16  cap16_1
timestamp 1667684462
transform 1 0 29700 0 1 6500
box 0 0 1450 6200
use cap16  cap16_2
timestamp 1667684462
transform 1 0 29700 0 -1 4900
box 0 0 1450 6200
use cap16  cap16_3
timestamp 1667684462
transform 1 0 24100 0 -1 4900
box 0 0 1450 6200
use cap32  cap32_0
timestamp 1667684412
transform 1 0 20900 0 1 6500
box 0 0 3050 6200
use cap32  cap32_1
timestamp 1667684412
transform 1 0 26500 0 1 6500
box 0 0 3050 6200
use cap32  cap32_2
timestamp 1667684412
transform 1 0 26500 0 -1 4900
box 0 0 3050 6200
use cap32  cap32_3
timestamp 1667684412
transform 1 0 20900 0 -1 4900
box 0 0 3050 6200
use cap64  cap64_0
timestamp 1667684360
transform 1 0 14500 0 1 6500
box 0 0 6250 6200
use cap64  cap64_1
timestamp 1667684360
transform 1 0 -4700 0 1 6500
box 0 0 6250 6200
use cap64  cap64_2
timestamp 1667684360
transform 1 0 14500 0 -1 4900
box 0 0 6250 6200
use cap64  cap64_3
timestamp 1667684360
transform 1 0 -4700 0 -1 4900
box 0 0 6250 6200
use cap128  cap128_0
timestamp 1667663783
transform 1 0 -17500 0 1 6500
box 0 0 12650 6200
use cap128  cap128_1
timestamp 1667663783
transform 1 0 1700 0 1 6500
box 0 0 12650 6200
use cap128  cap128_2
timestamp 1667663783
transform 1 0 1700 0 -1 4900
box 0 0 12650 6200
use cap128  cap128_3
timestamp 1667663783
transform 1 0 -17500 0 -1 4900
box 0 0 12650 6200
<< labels >>
rlabel metal4 43550 4100 43600 4300 1 sw_sp_n9
port 1 n
rlabel metal4 37150 4100 37200 4300 1 sw_sp_n8
port 2 n
rlabel metal4 35550 4100 36400 4250 1 sw_sp_n7
port 3 n
rlabel metal4 32350 4100 34800 4250 1 sw_sp_n6
port 4 n
rlabel metal4 25950 -1500 26000 -1100 1 sw_sp_n5
port 5 n
rlabel metal4 24350 -1500 25200 -1350 1 sw_sp_n4
port 6 n
rlabel metal4 21150 -1500 23600 -1350 1 sw_sp_n3
port 7 n
rlabel metal4 -4450 -1500 1200 -1350 1 sw_sp_n2
port 8 n
rlabel metal4 -17250 -1500 -5200 -1350 1 sw_sp_n1
port 9 n
rlabel metal4 -16910 6250 43950 6450 1 Vin_p
port 10 n
rlabel metal4 -16910 4950 43950 5150 1 Vin_n
port 11 n
rlabel metal4 43550 7100 43600 7300 1 sw_sp_p9
port 12 n
rlabel metal4 37150 7100 37200 7300 1 sw_sp_p8
port 13 n
rlabel metal4 35550 7150 36400 7300 1 sw_sp_p7
port 14 n
rlabel metal4 32350 7150 34800 7300 1 sw_sp_p6
port 15 n
rlabel metal4 25950 12500 26000 12900 1 sw_sp_p5
port 16 n
rlabel metal4 24350 12750 25200 12900 1 sw_sp_p4
port 17 n
rlabel metal4 21150 12750 23600 12900 1 sw_sp_p3
port 18 n
rlabel metal4 -4450 12750 1200 12900 1 sw_sp_p2
port 19 n
rlabel metal4 -17250 12750 -5200 12900 1 sw_sp_p1
port 20 n
rlabel metal4 42750 7100 42800 7300 1 sw_p8
port 21 n
rlabel metal4 41150 7150 42000 7300 1 sw_p7
port 22 n
rlabel metal4 37950 7150 40400 7300 1 sw_p6
port 23 n
rlabel metal4 31550 12500 31600 12900 1 sw_p5
port 24 n
rlabel metal4 29950 12750 30800 12900 1 sw_p4
port 25 n
rlabel metal4 26750 12750 29200 12900 1 sw_p3
port 26 n
rlabel metal4 14750 12750 20400 12900 1 sw_p2
port 27 n
rlabel metal4 1950 12750 14000 12900 1 sw_p1
port 28 n
rlabel metal4 42750 4100 42800 4300 1 sw_n8
port 29 n
rlabel metal4 41150 4100 42000 4250 1 sw_n7
port 30 n
rlabel metal4 37950 4100 40400 4250 1 sw_n6
port 31 n
rlabel metal4 31550 -1500 31600 -1100 1 sw_n5
port 32 n
rlabel metal4 29950 -1500 30800 -1350 1 sw_n4
port 33 n
rlabel metal4 26750 -1500 29200 -1350 1 sw_n3
port 34 n
rlabel metal4 14750 -1500 20400 -1350 1 sw_n2
port 35 n
rlabel metal4 1950 -1500 14000 -1350 1 sw_n1
port 36 n
<< end >>
