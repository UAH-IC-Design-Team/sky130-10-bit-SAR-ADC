magic
tech sky130A
magscale 1 2
timestamp 1666924247
<< nwell >>
rect -451 -269 449 221
<< pmos >>
rect -351 -161 -321 161
rect -255 -161 -225 161
rect -159 -161 -129 161
rect -63 -161 -33 161
rect 33 -161 63 161
rect 129 -161 159 161
rect 225 -161 255 161
rect 321 -161 351 161
<< pdiff >>
rect -413 149 -351 161
rect -413 -149 -401 149
rect -367 -149 -351 149
rect -413 -161 -351 -149
rect -321 149 -255 161
rect -321 -149 -305 149
rect -271 -149 -255 149
rect -321 -161 -255 -149
rect -225 149 -159 161
rect -225 -149 -209 149
rect -175 -149 -159 149
rect -225 -161 -159 -149
rect -129 149 -63 161
rect -129 -149 -113 149
rect -79 -149 -63 149
rect -129 -161 -63 -149
rect -33 149 33 161
rect -33 -149 -17 149
rect 17 -149 33 149
rect -33 -161 33 -149
rect 63 149 129 161
rect 63 -149 79 149
rect 113 -149 129 149
rect 63 -161 129 -149
rect 159 149 225 161
rect 159 -149 175 149
rect 209 -149 225 149
rect 159 -161 225 -149
rect 255 149 321 161
rect 255 -149 271 149
rect 305 -149 321 149
rect 255 -161 321 -149
rect 351 149 413 161
rect 351 -149 367 149
rect 401 -149 413 149
rect 351 -161 413 -149
<< pdiffc >>
rect -401 -149 -367 149
rect -305 -149 -271 149
rect -209 -149 -175 149
rect -113 -149 -79 149
rect -17 -149 17 149
rect 79 -149 113 149
rect 175 -149 209 149
rect 271 -149 305 149
rect 367 -149 401 149
<< poly >>
rect -351 161 -321 191
rect -255 161 -225 191
rect -159 161 -129 191
rect -63 161 -33 191
rect 33 161 63 191
rect 129 161 159 191
rect 225 161 255 191
rect 321 161 351 191
rect -351 -192 -321 -161
rect -255 -192 -225 -161
rect -159 -192 -129 -161
rect -63 -192 -33 -161
rect 33 -192 63 -161
rect 129 -192 159 -161
rect 225 -192 255 -161
rect 321 -192 351 -161
rect -377 -208 383 -192
rect -377 -242 -353 -208
rect -319 -242 -252 -208
rect -218 -242 -161 -208
rect -127 -242 -62 -208
rect -28 -242 31 -208
rect 65 -242 128 -208
rect 162 -242 223 -208
rect 257 -242 318 -208
rect 352 -242 383 -208
rect -377 -258 383 -242
<< polycont >>
rect -353 -242 -319 -208
rect -252 -242 -218 -208
rect -161 -242 -127 -208
rect -62 -242 -28 -208
rect 31 -242 65 -208
rect 128 -242 162 -208
rect 223 -242 257 -208
rect 318 -242 352 -208
<< locali >>
rect -401 149 -367 165
rect -401 -165 -367 -149
rect -305 149 -271 165
rect -305 -165 -271 -149
rect -209 149 -175 165
rect -209 -165 -175 -149
rect -113 149 -79 165
rect -113 -165 -79 -149
rect -17 149 17 165
rect -17 -165 17 -149
rect 79 149 113 165
rect 79 -165 113 -149
rect 175 149 209 165
rect 175 -165 209 -149
rect 271 149 305 165
rect 271 -165 305 -149
rect 367 149 401 165
rect 367 -165 401 -149
rect -377 -242 -353 -208
rect -319 -242 -252 -208
rect -218 -242 -161 -208
rect -127 -242 -62 -208
rect -28 -242 31 -208
rect 65 -242 128 -208
rect 162 -242 223 -208
rect 257 -242 318 -208
rect 352 -242 383 -208
<< viali >>
rect -401 28 -367 132
rect -305 -132 -271 -28
rect -209 28 -175 132
rect -113 -132 -79 -28
rect -17 28 17 132
rect 79 -132 113 -28
rect 175 28 209 132
rect 271 -132 305 -28
rect 367 28 401 132
rect -353 -242 -319 -208
rect -252 -242 -218 -208
rect -161 -242 -127 -208
rect -62 -242 -28 -208
rect 31 -242 65 -208
rect 128 -242 162 -208
rect 223 -242 257 -208
rect 318 -242 352 -208
<< metal1 >>
rect -407 132 -361 144
rect -407 28 -401 132
rect -367 28 -361 132
rect -407 16 -361 28
rect -215 132 -169 144
rect -215 28 -209 132
rect -175 28 -169 132
rect -215 16 -169 28
rect -23 132 23 144
rect -23 28 -17 132
rect 17 28 23 132
rect -23 16 23 28
rect 169 132 215 144
rect 169 28 175 132
rect 209 28 215 132
rect 169 16 215 28
rect 361 132 407 144
rect 361 28 367 132
rect 401 28 407 132
rect 361 16 407 28
rect -311 -28 -265 -16
rect -311 -132 -305 -28
rect -271 -132 -265 -28
rect -311 -144 -265 -132
rect -119 -28 -73 -16
rect -119 -132 -113 -28
rect -79 -132 -73 -28
rect -119 -144 -73 -132
rect 73 -28 119 -16
rect 73 -132 79 -28
rect 113 -132 119 -28
rect 73 -144 119 -132
rect 265 -28 311 -16
rect 265 -132 271 -28
rect 305 -132 311 -28
rect 265 -144 311 -132
rect -377 -208 383 -202
rect -377 -242 -353 -208
rect -319 -242 -252 -208
rect -218 -242 -161 -208
rect -127 -242 -62 -208
rect -28 -242 31 -208
rect 65 -242 128 -208
rect 162 -242 223 -208
rect 257 -242 318 -208
rect 352 -242 383 -208
rect -377 -248 383 -242
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc +35 viadrn -35 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
