magic
tech sky130A
magscale 1 2
timestamp 1666551745
<< nwell >>
rect -20 1080 1980 2060
<< psubdiff >>
rect 360 910 420 934
rect 360 746 420 770
rect 580 680 640 704
rect 580 516 640 540
rect 726 470 750 540
rect 940 470 964 540
rect 1100 440 1160 464
rect 1100 276 1160 300
rect 1226 90 1250 150
rect 1440 90 1464 150
<< nsubdiff >>
rect 1090 1920 1120 1980
rect 1210 1920 1240 1980
rect 1090 1780 1120 1840
rect 1210 1780 1240 1840
rect 1090 1640 1120 1700
rect 1210 1640 1240 1700
rect 600 1450 630 1510
rect 720 1450 750 1510
rect 170 1380 200 1440
rect 290 1380 320 1440
<< psubdiffcont >>
rect 360 770 420 910
rect 580 540 640 680
rect 750 470 940 540
rect 1100 300 1160 440
rect 1250 90 1440 150
<< nsubdiffcont >>
rect 1120 1920 1210 1980
rect 1120 1780 1210 1840
rect 1120 1640 1210 1700
rect 630 1450 720 1510
rect 200 1380 290 1440
<< locali >>
rect 1100 1920 1120 1980
rect 1210 1920 1230 1980
rect 1100 1780 1120 1840
rect 1210 1780 1230 1840
rect 1100 1640 1120 1700
rect 1210 1640 1230 1700
rect 610 1450 630 1510
rect 720 1450 740 1510
rect 180 1380 200 1440
rect 290 1380 310 1440
rect 360 910 420 926
rect 360 760 370 770
rect 410 760 420 770
rect 360 754 420 760
rect 580 680 640 696
rect 580 524 640 540
rect 734 470 750 540
rect 940 470 956 540
rect 1100 440 1160 456
rect 1100 284 1160 300
rect 1234 90 1250 150
rect 1440 90 1456 150
<< viali >>
rect 1120 1920 1210 1980
rect 1120 1780 1210 1840
rect 1120 1640 1210 1700
rect 630 1450 720 1510
rect 200 1380 290 1440
rect 370 770 410 890
rect 370 760 410 770
rect 590 540 630 670
rect 760 480 930 530
rect 1110 300 1150 440
rect 1250 100 1430 140
<< metal1 >>
rect 1100 1980 1750 2030
rect 1090 1920 1120 1980
rect 1210 1940 1750 1980
rect 1210 1920 1240 1940
rect 1100 1840 1230 1920
rect 1090 1780 1120 1840
rect 1210 1780 1240 1840
rect 1100 1700 1230 1780
rect 1090 1640 1120 1700
rect 1210 1640 1240 1700
rect 620 1580 1230 1640
rect 620 1510 730 1580
rect 600 1450 630 1510
rect 720 1450 750 1510
rect 180 1440 730 1450
rect 180 1380 200 1440
rect 290 1380 730 1440
rect -20 900 40 1220
rect 180 1210 310 1380
rect 90 1080 250 1170
rect 480 1080 540 1340
rect 620 1220 730 1380
rect 760 1090 900 1360
rect 1000 1090 1060 1540
rect 1110 1220 1230 1580
rect 1270 1090 1410 1550
rect 1520 1090 1580 1900
rect 1630 1220 1750 1940
rect 1790 1110 1930 1940
rect 90 1020 540 1080
rect 90 960 250 1020
rect 70 890 420 910
rect 70 860 370 890
rect 360 760 370 860
rect 410 760 420 890
rect 480 800 540 1020
rect 680 1030 1060 1090
rect 580 760 640 910
rect 680 760 740 1030
rect 360 710 640 760
rect 580 670 640 710
rect 580 540 590 670
rect 630 540 640 670
rect 1000 580 1060 1030
rect 1200 1030 1580 1090
rect 1100 540 1160 900
rect 1200 560 1270 1030
rect 580 530 1160 540
rect 580 480 760 530
rect 930 480 1160 530
rect 580 470 1160 480
rect 1100 440 1160 470
rect 1100 300 1110 440
rect 1150 300 1160 440
rect 1100 150 1160 300
rect 1520 200 1580 1030
rect 1720 1010 1980 1110
rect 1620 150 1680 910
rect 1720 180 1810 1010
rect 1100 140 1680 150
rect 1100 100 1250 140
rect 1430 100 1680 140
rect 1100 90 1680 100
use sky130_fd_pr__nfet_01v8_9CGS2F  XM1
timestamp 1666487809
transform 0 1 128 -1 0 933
box -73 -148 73 148
use sky130_fd_pr__pfet_01v8_46WN3R  XM2
timestamp 1666487809
transform 0 1 209 1 0 1189
box -109 -229 109 263
use sky130_fd_pr__nfet_01v8_5XXJZ8  XM3
timestamp 1666487809
transform 0 1 659 -1 0 885
box -125 -179 125 121
use sky130_fd_pr__pfet_01v8_CBMBZG  XM4
timestamp 1666490112
transform 0 1 745 -1 0 1241
box -169 -265 161 205
use sky130_fd_pr__nfet_01v8_ZDVJZL  XM5
timestamp 1666489008
transform 0 1 1179 -1 0 781
box -221 -179 221 121
use sky130_fd_pr__pfet_01v8_CBDHKH  XM6
timestamp 1666490340
transform 0 1 1255 -1 0 1337
box -263 -265 257 205
use sky130_fd_pr__nfet_01v8_MRXJZU  XM7
timestamp 1666489318
transform 0 1 1699 -1 0 593
box -413 -179 413 121
use sky130_fd_pr__pfet_01v8_CBVRKH  XM8
timestamp 1666490724
transform 0 1 1775 -1 0 1529
box -451 -265 449 205
<< labels >>
rlabel metal1 1210 1940 1750 2030 1 VDD
port 1 n
rlabel metal1 -20 900 40 1220 1 Vin
port 2 n
rlabel metal1 1720 1010 1980 1110 1 Vout
port 3 n
rlabel metal1 1100 90 1680 150 1 VSS
port 4 n
<< end >>
