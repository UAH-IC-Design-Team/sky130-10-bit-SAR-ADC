magic
tech sky130A
magscale 1 2
timestamp 1666377729
<< error_p >>
rect -77 246 -19 252
rect 115 246 173 252
rect -77 212 -65 246
rect 115 212 127 246
rect -77 206 -19 212
rect 115 206 173 212
rect -173 -212 -115 -206
rect 19 -212 77 -206
rect -173 -246 -161 -212
rect 19 -246 31 -212
rect -173 -252 -115 -246
rect 19 -252 77 -246
<< nwell >>
rect -161 227 257 265
rect -257 -227 257 227
rect -257 -265 161 -227
<< pmos >>
rect -159 -165 -129 165
rect -63 -165 -33 165
rect 33 -165 63 165
rect 129 -165 159 165
<< pdiff >>
rect -221 153 -159 165
rect -221 -153 -209 153
rect -175 -153 -159 153
rect -221 -165 -159 -153
rect -129 153 -63 165
rect -129 -153 -113 153
rect -79 -153 -63 153
rect -129 -165 -63 -153
rect -33 153 33 165
rect -33 -153 -17 153
rect 17 -153 33 153
rect -33 -165 33 -153
rect 63 153 129 165
rect 63 -153 79 153
rect 113 -153 129 153
rect 63 -165 129 -153
rect 159 153 221 165
rect 159 -153 175 153
rect 209 -153 221 153
rect 159 -165 221 -153
<< pdiffc >>
rect -209 -153 -175 153
rect -113 -153 -79 153
rect -17 -153 17 153
rect 79 -153 113 153
rect 175 -153 209 153
<< poly >>
rect -81 246 -15 262
rect -81 212 -65 246
rect -31 212 -15 246
rect -81 196 -15 212
rect 111 246 177 262
rect 111 212 127 246
rect 161 212 177 246
rect 111 196 177 212
rect -159 165 -129 191
rect -63 165 -33 196
rect 33 165 63 191
rect 129 165 159 196
rect -159 -196 -129 -165
rect -63 -191 -33 -165
rect 33 -196 63 -165
rect 129 -191 159 -165
rect -177 -212 -111 -196
rect -177 -246 -161 -212
rect -127 -246 -111 -212
rect -177 -262 -111 -246
rect 15 -212 81 -196
rect 15 -246 31 -212
rect 65 -246 81 -212
rect 15 -262 81 -246
<< polycont >>
rect -65 212 -31 246
rect 127 212 161 246
rect -161 -246 -127 -212
rect 31 -246 65 -212
<< locali >>
rect -81 212 -65 246
rect -31 212 -15 246
rect 111 212 127 246
rect 161 212 177 246
rect -209 153 -175 169
rect -209 -169 -175 -153
rect -113 153 -79 169
rect -113 -169 -79 -153
rect -17 153 17 169
rect -17 -169 17 -153
rect 79 153 113 169
rect 79 -169 113 -153
rect 175 153 209 169
rect 175 -169 209 -153
rect -177 -246 -161 -212
rect -127 -246 -111 -212
rect 15 -246 31 -212
rect 65 -246 81 -212
<< viali >>
rect -65 212 -31 246
rect 127 212 161 246
rect -209 -153 -175 153
rect -113 -136 -79 -29
rect -17 -153 17 153
rect 79 -136 113 -29
rect 175 -153 209 153
rect -161 -246 -127 -212
rect 31 -246 65 -212
<< metal1 >>
rect -77 246 -19 252
rect -77 212 -65 246
rect -31 212 -19 246
rect -77 206 -19 212
rect 115 246 173 252
rect 115 212 127 246
rect 161 212 173 246
rect 115 206 173 212
rect -215 153 -169 165
rect -215 -153 -209 153
rect -175 -153 -169 153
rect -23 153 23 165
rect -119 -29 -73 -17
rect -119 -136 -113 -29
rect -79 -136 -73 -29
rect -119 -148 -73 -136
rect -215 -165 -169 -153
rect -23 -153 -17 153
rect 17 -153 23 153
rect 169 153 215 165
rect 73 -29 119 -17
rect 73 -136 79 -29
rect 113 -136 119 -29
rect 73 -148 119 -136
rect -23 -165 23 -153
rect 169 -153 175 153
rect 209 -153 215 153
rect 169 -165 215 -153
rect -173 -212 -115 -206
rect -173 -246 -161 -212
rect -127 -246 -115 -212
rect -173 -252 -115 -246
rect 19 -212 77 -206
rect 19 -246 31 -212
rect 65 -246 77 -212
rect 19 -252 77 -246
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc +35 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
