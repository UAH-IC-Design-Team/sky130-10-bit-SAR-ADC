magic
tech sky130A
magscale 1 2
timestamp 1666650150
<< error_p >>
rect -125 181 -67 187
rect 67 181 125 187
rect -125 147 -113 181
rect 67 147 79 181
rect -125 141 -67 147
rect 67 141 125 147
rect -221 -147 -163 -141
rect -29 -147 29 -141
rect 163 -147 221 -141
rect -221 -181 -209 -147
rect -29 -181 -17 -147
rect 163 -181 175 -147
rect -221 -187 -163 -181
rect -29 -187 29 -181
rect 163 -187 221 -181
<< nwell >>
rect -407 -319 407 319
<< pmos >>
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
<< pdiff >>
rect -269 88 -207 100
rect -269 -88 -257 88
rect -223 -88 -207 88
rect -269 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 269 100
rect 207 -88 223 88
rect 257 -88 269 88
rect 207 -100 269 -88
<< pdiffc >>
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
<< nsubdiff >>
rect -371 249 -275 283
rect 275 249 371 283
rect -371 187 -337 249
rect 337 187 371 249
rect -371 -249 -337 -187
rect 337 -249 371 -187
rect -371 -283 -275 -249
rect 275 -283 371 -249
<< nsubdiffcont >>
rect -275 249 275 283
rect -371 -187 -337 187
rect 337 -187 371 187
rect -275 -283 275 -249
<< poly >>
rect -129 181 -63 197
rect -129 147 -113 181
rect -79 147 -63 181
rect -129 131 -63 147
rect 63 181 129 197
rect 63 147 79 181
rect 113 147 129 181
rect 63 131 129 147
rect -207 100 -177 126
rect -111 100 -81 131
rect -15 100 15 126
rect 81 100 111 131
rect 177 100 207 126
rect -207 -131 -177 -100
rect -111 -126 -81 -100
rect -15 -131 15 -100
rect 81 -126 111 -100
rect 177 -131 207 -100
rect -225 -147 -159 -131
rect -225 -181 -209 -147
rect -175 -181 -159 -147
rect -225 -197 -159 -181
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
rect 159 -147 225 -131
rect 159 -181 175 -147
rect 209 -181 225 -147
rect 159 -197 225 -181
<< polycont >>
rect -113 147 -79 181
rect 79 147 113 181
rect -209 -181 -175 -147
rect -17 -181 17 -147
rect 175 -181 209 -147
<< locali >>
rect -371 249 -275 283
rect 275 249 371 283
rect -371 187 -337 249
rect 337 187 371 249
rect -129 147 -113 181
rect -79 147 -63 181
rect 63 147 79 181
rect 113 147 129 181
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect -225 -181 -209 -147
rect -175 -181 -159 -147
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect 159 -181 175 -147
rect 209 -181 225 -147
rect -371 -249 -337 -187
rect 337 -249 371 -187
rect -371 -283 -275 -249
rect 275 -283 371 -249
<< viali >>
rect -113 147 -79 181
rect 79 147 113 181
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect -209 -181 -175 -147
rect -17 -181 17 -147
rect 175 -181 209 -147
<< metal1 >>
rect -125 181 -67 187
rect -125 147 -113 181
rect -79 147 -67 181
rect -125 141 -67 147
rect 67 181 125 187
rect 67 147 79 181
rect 113 147 125 181
rect 67 141 125 147
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect -221 -147 -163 -141
rect -221 -181 -209 -147
rect -175 -181 -163 -147
rect -221 -187 -163 -181
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
rect 163 -147 221 -141
rect 163 -181 175 -147
rect 209 -181 221 -147
rect 163 -187 221 -181
<< properties >>
string FIXED_BBOX -354 -266 354 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
