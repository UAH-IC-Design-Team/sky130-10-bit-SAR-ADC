magic
tech sky130A
magscale 1 2
timestamp 1666918349
<< error_p >>
rect -29 1079 29 1085
rect -29 1045 -17 1079
rect -29 1039 29 1045
rect -29 629 29 635
rect -29 595 -17 629
rect -29 589 29 595
rect -29 521 29 527
rect -29 487 -17 521
rect -29 481 29 487
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -487 29 -481
rect -29 -521 -17 -487
rect -29 -527 29 -521
rect -29 -595 29 -589
rect -29 -629 -17 -595
rect -29 -635 29 -629
rect -29 -1045 29 -1039
rect -29 -1079 -17 -1045
rect -29 -1085 29 -1079
<< nwell >>
rect -211 -1217 211 1217
<< pmos >>
rect -15 676 15 998
rect -15 118 15 440
rect -15 -440 15 -118
rect -15 -998 15 -676
<< pdiff >>
rect -73 986 -15 998
rect -73 688 -61 986
rect -27 688 -15 986
rect -73 676 -15 688
rect 15 986 73 998
rect 15 688 27 986
rect 61 688 73 986
rect 15 676 73 688
rect -73 428 -15 440
rect -73 130 -61 428
rect -27 130 -15 428
rect -73 118 -15 130
rect 15 428 73 440
rect 15 130 27 428
rect 61 130 73 428
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -428 -61 -130
rect -27 -428 -15 -130
rect -73 -440 -15 -428
rect 15 -130 73 -118
rect 15 -428 27 -130
rect 61 -428 73 -130
rect 15 -440 73 -428
rect -73 -688 -15 -676
rect -73 -986 -61 -688
rect -27 -986 -15 -688
rect -73 -998 -15 -986
rect 15 -688 73 -676
rect 15 -986 27 -688
rect 61 -986 73 -688
rect 15 -998 73 -986
<< pdiffc >>
rect -61 688 -27 986
rect 27 688 61 986
rect -61 130 -27 428
rect 27 130 61 428
rect -61 -428 -27 -130
rect 27 -428 61 -130
rect -61 -986 -27 -688
rect 27 -986 61 -688
<< nsubdiff >>
rect -175 1147 -79 1181
rect 79 1147 175 1181
rect -175 1085 -141 1147
rect 141 1085 175 1147
rect -175 -1147 -141 -1085
rect 141 -1147 175 -1085
rect -175 -1181 -79 -1147
rect 79 -1181 175 -1147
<< nsubdiffcont >>
rect -79 1147 79 1181
rect -175 -1085 -141 1085
rect 141 -1085 175 1085
rect -79 -1181 79 -1147
<< poly >>
rect -33 1079 33 1095
rect -33 1045 -17 1079
rect 17 1045 33 1079
rect -33 1029 33 1045
rect -15 998 15 1029
rect -15 645 15 676
rect -33 629 33 645
rect -33 595 -17 629
rect 17 595 33 629
rect -33 579 33 595
rect -33 521 33 537
rect -33 487 -17 521
rect 17 487 33 521
rect -33 471 33 487
rect -15 440 15 471
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -471 15 -440
rect -33 -487 33 -471
rect -33 -521 -17 -487
rect 17 -521 33 -487
rect -33 -537 33 -521
rect -33 -595 33 -579
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -33 -645 33 -629
rect -15 -676 15 -645
rect -15 -1029 15 -998
rect -33 -1045 33 -1029
rect -33 -1079 -17 -1045
rect 17 -1079 33 -1045
rect -33 -1095 33 -1079
<< polycont >>
rect -17 1045 17 1079
rect -17 595 17 629
rect -17 487 17 521
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -521 17 -487
rect -17 -629 17 -595
rect -17 -1079 17 -1045
<< locali >>
rect -175 1147 -79 1181
rect 79 1147 175 1181
rect -175 1085 -141 1147
rect 141 1085 175 1147
rect -33 1045 -17 1079
rect 17 1045 33 1079
rect -61 986 -27 1002
rect -61 672 -27 688
rect 27 986 61 1002
rect 27 672 61 688
rect -33 595 -17 629
rect 17 595 33 629
rect -33 487 -17 521
rect 17 487 33 521
rect -61 428 -27 444
rect -61 114 -27 130
rect 27 428 61 444
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -444 -27 -428
rect 27 -130 61 -114
rect 27 -444 61 -428
rect -33 -521 -17 -487
rect 17 -521 33 -487
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -61 -688 -27 -672
rect -61 -1002 -27 -986
rect 27 -688 61 -672
rect 27 -1002 61 -986
rect -33 -1079 -17 -1045
rect 17 -1079 33 -1045
rect -175 -1147 -141 -1085
rect 141 -1147 175 -1085
rect -175 -1181 -79 -1147
rect 79 -1181 175 -1147
<< viali >>
rect -17 1045 17 1079
rect -61 688 -27 986
rect 27 688 61 986
rect -17 595 17 629
rect -17 487 17 521
rect -61 130 -27 428
rect 27 130 61 428
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -428 -27 -130
rect 27 -428 61 -130
rect -17 -521 17 -487
rect -17 -629 17 -595
rect -61 -986 -27 -688
rect 27 -986 61 -688
rect -17 -1079 17 -1045
<< metal1 >>
rect -29 1079 29 1085
rect -29 1045 -17 1079
rect 17 1045 29 1079
rect -29 1039 29 1045
rect -67 986 -21 998
rect -67 688 -61 986
rect -27 688 -21 986
rect -67 676 -21 688
rect 21 986 67 998
rect 21 688 27 986
rect 61 688 67 986
rect 21 676 67 688
rect -29 629 29 635
rect -29 595 -17 629
rect 17 595 29 629
rect -29 589 29 595
rect -29 521 29 527
rect -29 487 -17 521
rect 17 487 29 521
rect -29 481 29 487
rect -67 428 -21 440
rect -67 130 -61 428
rect -27 130 -21 428
rect -67 118 -21 130
rect 21 428 67 440
rect 21 130 27 428
rect 61 130 67 428
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -428 -61 -130
rect -27 -428 -21 -130
rect -67 -440 -21 -428
rect 21 -130 67 -118
rect 21 -428 27 -130
rect 61 -428 67 -130
rect 21 -440 67 -428
rect -29 -487 29 -481
rect -29 -521 -17 -487
rect 17 -521 29 -487
rect -29 -527 29 -521
rect -29 -595 29 -589
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -635 29 -629
rect -67 -688 -21 -676
rect -67 -986 -61 -688
rect -27 -986 -21 -688
rect -67 -998 -21 -986
rect 21 -688 67 -676
rect 21 -986 27 -688
rect 61 -986 67 -688
rect 21 -998 67 -986
rect -29 -1045 29 -1039
rect -29 -1079 -17 -1045
rect 17 -1079 29 -1045
rect -29 -1085 29 -1079
<< properties >>
string FIXED_BBOX -158 -1164 158 1164
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
