magic
tech sky130A
magscale 1 2
timestamp 1667686553
<< metal1 >>
rect -33560 12220 -33140 12240
rect -33560 12080 -33540 12220
rect -33160 12080 -33140 12220
rect -33560 12060 -33140 12080
<< via1 >>
rect -33540 12080 -33160 12220
<< metal2 >>
rect -33560 12220 -33140 12240
rect -33560 12080 -33540 12220
rect -33160 12080 -33140 12220
rect -33560 12060 -33140 12080
<< via2 >>
rect -33540 12080 -33160 12220
<< metal3 >>
rect -33340 12880 -32400 12900
rect -33340 12740 -33320 12880
rect -33040 12740 -32680 12880
rect -32420 12740 -32400 12880
rect -33340 12660 -32400 12740
rect -33340 12520 -33320 12660
rect -33040 12520 -32680 12660
rect -32420 12520 -32400 12660
rect -33340 12500 -32400 12520
rect -31740 12880 -30800 12900
rect -31740 12740 -31720 12880
rect -31440 12740 -31080 12880
rect -30820 12740 -30800 12880
rect -31740 12660 -30800 12740
rect -31740 12520 -31720 12660
rect -31440 12520 -31080 12660
rect -30820 12520 -30800 12660
rect -31740 12500 -30800 12520
rect -30140 12880 -29200 12900
rect -30140 12740 -30120 12880
rect -29840 12740 -29480 12880
rect -29220 12740 -29200 12880
rect -30140 12660 -29200 12740
rect -30140 12520 -30120 12660
rect -29840 12520 -29480 12660
rect -29220 12520 -29200 12660
rect -30140 12500 -29200 12520
rect -28540 12880 -27600 12900
rect -28540 12740 -28520 12880
rect -28240 12740 -27880 12880
rect -27620 12740 -27600 12880
rect -28540 12660 -27600 12740
rect -28540 12520 -28520 12660
rect -28240 12520 -27880 12660
rect -27620 12520 -27600 12660
rect -28540 12500 -27600 12520
rect -26940 12880 -26000 12900
rect -26940 12740 -26920 12880
rect -26640 12740 -26280 12880
rect -26020 12740 -26000 12880
rect -26940 12660 -26000 12740
rect -26940 12520 -26920 12660
rect -26640 12520 -26280 12660
rect -26020 12520 -26000 12660
rect -26940 12500 -26000 12520
rect -25340 12880 -24400 12900
rect -25340 12740 -25320 12880
rect -25040 12740 -24680 12880
rect -24420 12740 -24400 12880
rect -25340 12660 -24400 12740
rect -25340 12520 -25320 12660
rect -25040 12520 -24680 12660
rect -24420 12520 -24400 12660
rect -25340 12500 -24400 12520
rect -23740 12880 -22800 12900
rect -23740 12740 -23720 12880
rect -23440 12740 -23080 12880
rect -22820 12740 -22800 12880
rect -23740 12660 -22800 12740
rect -23740 12520 -23720 12660
rect -23440 12520 -23080 12660
rect -22820 12520 -22800 12660
rect -23740 12500 -22800 12520
rect -22140 12880 -21200 12900
rect -22140 12740 -22120 12880
rect -21840 12740 -21480 12880
rect -21220 12740 -21200 12880
rect -22140 12660 -21200 12740
rect -22140 12520 -22120 12660
rect -21840 12520 -21480 12660
rect -21220 12520 -21200 12660
rect -22140 12500 -21200 12520
rect -20540 12880 -19600 12900
rect -20540 12740 -20520 12880
rect -20240 12740 -19880 12880
rect -19620 12740 -19600 12880
rect -20540 12660 -19600 12740
rect -20540 12520 -20520 12660
rect -20240 12520 -19880 12660
rect -19620 12520 -19600 12660
rect -20540 12500 -19600 12520
rect -18940 12880 -18000 12900
rect -18940 12740 -18920 12880
rect -18640 12740 -18280 12880
rect -18020 12740 -18000 12880
rect -18940 12660 -18000 12740
rect -18940 12520 -18920 12660
rect -18640 12520 -18280 12660
rect -18020 12520 -18000 12660
rect -18940 12500 -18000 12520
rect -17340 12880 -16400 12900
rect -17340 12740 -17320 12880
rect -17040 12740 -16680 12880
rect -16420 12740 -16400 12880
rect -17340 12660 -16400 12740
rect -17340 12520 -17320 12660
rect -17040 12520 -16680 12660
rect -16420 12520 -16400 12660
rect -17340 12500 -16400 12520
rect -15740 12880 -14800 12900
rect -15740 12740 -15720 12880
rect -15440 12740 -15080 12880
rect -14820 12740 -14800 12880
rect -15740 12660 -14800 12740
rect -15740 12520 -15720 12660
rect -15440 12520 -15080 12660
rect -14820 12520 -14800 12660
rect -15740 12500 -14800 12520
rect -14140 12880 -13200 12900
rect -14140 12740 -14120 12880
rect -13840 12740 -13480 12880
rect -13220 12740 -13200 12880
rect -14140 12660 -13200 12740
rect -14140 12520 -14120 12660
rect -13840 12520 -13480 12660
rect -13220 12520 -13200 12660
rect -14140 12500 -13200 12520
rect -12540 12880 -11600 12900
rect -12540 12740 -12520 12880
rect -12240 12740 -11880 12880
rect -11620 12740 -11600 12880
rect -12540 12660 -11600 12740
rect -12540 12520 -12520 12660
rect -12240 12520 -11880 12660
rect -11620 12520 -11600 12660
rect -12540 12500 -11600 12520
rect -10940 12880 -10000 12900
rect -10940 12740 -10920 12880
rect -10640 12740 -10280 12880
rect -10020 12740 -10000 12880
rect -10940 12660 -10000 12740
rect -10940 12520 -10920 12660
rect -10640 12520 -10280 12660
rect -10020 12520 -10000 12660
rect -10940 12500 -10000 12520
rect -9340 12880 -8400 12900
rect -9340 12740 -9320 12880
rect -9040 12740 -8680 12880
rect -8420 12740 -8400 12880
rect -9340 12660 -8400 12740
rect -9340 12520 -9320 12660
rect -9040 12520 -8680 12660
rect -8420 12520 -8400 12660
rect -9340 12500 -8400 12520
rect -7740 12880 -6800 12900
rect -7740 12740 -7720 12880
rect -7440 12740 -7080 12880
rect -6820 12740 -6800 12880
rect -7740 12660 -6800 12740
rect -7740 12520 -7720 12660
rect -7440 12520 -7080 12660
rect -6820 12520 -6800 12660
rect -7740 12500 -6800 12520
rect -6140 12880 -5200 12900
rect -6140 12740 -6120 12880
rect -5840 12740 -5480 12880
rect -5220 12740 -5200 12880
rect -6140 12660 -5200 12740
rect -6140 12520 -6120 12660
rect -5840 12520 -5480 12660
rect -5220 12520 -5200 12660
rect -6140 12500 -5200 12520
rect -4540 12880 -3600 12900
rect -4540 12740 -4520 12880
rect -4240 12740 -3880 12880
rect -3620 12740 -3600 12880
rect -4540 12660 -3600 12740
rect -4540 12520 -4520 12660
rect -4240 12520 -3880 12660
rect -3620 12520 -3600 12660
rect -4540 12500 -3600 12520
rect -2940 12880 -2000 12900
rect -2940 12740 -2920 12880
rect -2640 12740 -2280 12880
rect -2020 12740 -2000 12880
rect -2940 12660 -2000 12740
rect -2940 12520 -2920 12660
rect -2640 12520 -2280 12660
rect -2020 12520 -2000 12660
rect -2940 12500 -2000 12520
rect -1340 12880 -400 12900
rect -1340 12740 -1320 12880
rect -1040 12740 -680 12880
rect -420 12740 -400 12880
rect -1340 12660 -400 12740
rect -1340 12520 -1320 12660
rect -1040 12520 -680 12660
rect -420 12520 -400 12660
rect -1340 12500 -400 12520
rect 260 12880 1200 12900
rect 260 12740 280 12880
rect 560 12740 920 12880
rect 1180 12740 1200 12880
rect 260 12660 1200 12740
rect 260 12520 280 12660
rect 560 12520 920 12660
rect 1180 12520 1200 12660
rect 260 12500 1200 12520
rect 1860 12880 2800 12900
rect 1860 12740 1880 12880
rect 2160 12740 2520 12880
rect 2780 12740 2800 12880
rect 1860 12660 2800 12740
rect 1860 12520 1880 12660
rect 2160 12520 2520 12660
rect 2780 12520 2800 12660
rect 1860 12500 2800 12520
rect 3460 12880 4400 12900
rect 3460 12740 3480 12880
rect 3760 12740 4120 12880
rect 4380 12740 4400 12880
rect 3460 12660 4400 12740
rect 3460 12520 3480 12660
rect 3760 12520 4120 12660
rect 4380 12520 4400 12660
rect 3460 12500 4400 12520
rect 5060 12880 6000 12900
rect 5060 12740 5080 12880
rect 5360 12740 5720 12880
rect 5980 12740 6000 12880
rect 5060 12660 6000 12740
rect 5060 12520 5080 12660
rect 5360 12520 5720 12660
rect 5980 12520 6000 12660
rect 5060 12500 6000 12520
rect 6660 12880 7600 12900
rect 6660 12740 6680 12880
rect 6960 12740 7320 12880
rect 7580 12740 7600 12880
rect 6660 12660 7600 12740
rect 6660 12520 6680 12660
rect 6960 12520 7320 12660
rect 7580 12520 7600 12660
rect 6660 12500 7600 12520
rect 8260 12880 9200 12900
rect 8260 12740 8280 12880
rect 8560 12740 8920 12880
rect 9180 12740 9200 12880
rect 8260 12660 9200 12740
rect 8260 12520 8280 12660
rect 8560 12520 8920 12660
rect 9180 12520 9200 12660
rect 8260 12500 9200 12520
rect 9860 12880 10800 12900
rect 9860 12740 9880 12880
rect 10160 12740 10520 12880
rect 10780 12740 10800 12880
rect 9860 12660 10800 12740
rect 9860 12520 9880 12660
rect 10160 12520 10520 12660
rect 10780 12520 10800 12660
rect 9860 12500 10800 12520
rect 11460 12880 12400 12900
rect 11460 12740 11480 12880
rect 11760 12740 12120 12880
rect 12380 12740 12400 12880
rect 11460 12660 12400 12740
rect 11460 12520 11480 12660
rect 11760 12520 12120 12660
rect 12380 12520 12400 12660
rect 11460 12500 12400 12520
rect 13060 12880 14000 12900
rect 13060 12740 13080 12880
rect 13360 12740 13720 12880
rect 13980 12740 14000 12880
rect 13060 12660 14000 12740
rect 13060 12520 13080 12660
rect 13360 12520 13720 12660
rect 13980 12520 14000 12660
rect 13060 12500 14000 12520
rect 14660 12880 15600 12900
rect 14660 12740 14680 12880
rect 14960 12740 15320 12880
rect 15580 12740 15600 12880
rect 14660 12660 15600 12740
rect 14660 12520 14680 12660
rect 14960 12520 15320 12660
rect 15580 12520 15600 12660
rect 14660 12500 15600 12520
rect 16260 12880 17200 12900
rect 16260 12740 16280 12880
rect 16560 12740 16920 12880
rect 17180 12740 17200 12880
rect 16260 12660 17200 12740
rect 16260 12520 16280 12660
rect 16560 12520 16920 12660
rect 17180 12520 17200 12660
rect 16260 12500 17200 12520
rect 17860 12880 18800 12900
rect 17860 12740 17880 12880
rect 18160 12740 18520 12880
rect 18780 12740 18800 12880
rect 17860 12660 18800 12740
rect 17860 12520 17880 12660
rect 18160 12520 18520 12660
rect 18780 12520 18800 12660
rect 17860 12500 18800 12520
rect 19460 12880 20400 12900
rect 19460 12740 19480 12880
rect 19760 12740 20120 12880
rect 20380 12740 20400 12880
rect 19460 12660 20400 12740
rect 19460 12520 19480 12660
rect 19760 12520 20120 12660
rect 20380 12520 20400 12660
rect 19460 12500 20400 12520
rect 21060 12880 22000 12900
rect 21060 12740 21080 12880
rect 21360 12740 21720 12880
rect 21980 12740 22000 12880
rect 21060 12660 22000 12740
rect 21060 12520 21080 12660
rect 21360 12520 21720 12660
rect 21980 12520 22000 12660
rect 21060 12500 22000 12520
rect 22660 12880 23600 12900
rect 22660 12740 22680 12880
rect 22960 12740 23320 12880
rect 23580 12740 23600 12880
rect 22660 12660 23600 12740
rect 22660 12520 22680 12660
rect 22960 12520 23320 12660
rect 23580 12520 23600 12660
rect 22660 12500 23600 12520
rect 24260 12880 25200 12900
rect 24260 12740 24280 12880
rect 24560 12740 24920 12880
rect 25180 12740 25200 12880
rect 24260 12660 25200 12740
rect 24260 12520 24280 12660
rect 24560 12520 24920 12660
rect 25180 12520 25200 12660
rect 24260 12500 25200 12520
rect 25860 12880 26800 12900
rect 25860 12740 25880 12880
rect 26160 12740 26520 12880
rect 26780 12740 26800 12880
rect 25860 12660 26800 12740
rect 25860 12520 25880 12660
rect 26160 12520 26520 12660
rect 26780 12520 26800 12660
rect 25860 12500 26800 12520
rect 27460 12880 28400 12900
rect 27460 12740 27480 12880
rect 27760 12740 28120 12880
rect 28380 12740 28400 12880
rect 27460 12660 28400 12740
rect 27460 12520 27480 12660
rect 27760 12520 28120 12660
rect 28380 12520 28400 12660
rect 27460 12500 28400 12520
rect 29060 12880 30000 12900
rect 29060 12740 29080 12880
rect 29360 12740 29720 12880
rect 29980 12740 30000 12880
rect 29060 12660 30000 12740
rect 29060 12520 29080 12660
rect 29360 12520 29720 12660
rect 29980 12520 30000 12660
rect 29060 12500 30000 12520
rect 30660 12880 31600 12900
rect 30660 12740 30680 12880
rect 30960 12740 31320 12880
rect 31580 12740 31600 12880
rect 30660 12660 31600 12740
rect 30660 12520 30680 12660
rect 30960 12520 31320 12660
rect 31580 12520 31600 12660
rect 30660 12500 31600 12520
rect 32260 12880 33200 12900
rect 32260 12740 32280 12880
rect 32560 12740 32920 12880
rect 33180 12740 33200 12880
rect 32260 12660 33200 12740
rect 32260 12520 32280 12660
rect 32560 12520 32920 12660
rect 33180 12520 33200 12660
rect 32260 12500 33200 12520
rect 33860 12880 34800 12900
rect 33860 12740 33880 12880
rect 34160 12740 34520 12880
rect 34780 12740 34800 12880
rect 33860 12660 34800 12740
rect 33860 12520 33880 12660
rect 34160 12520 34520 12660
rect 34780 12520 34800 12660
rect 33860 12500 34800 12520
rect 35460 12880 36400 12900
rect 35460 12740 35480 12880
rect 35760 12740 36120 12880
rect 36380 12740 36400 12880
rect 35460 12660 36400 12740
rect 35460 12520 35480 12660
rect 35760 12520 36120 12660
rect 36380 12520 36400 12660
rect 35460 12500 36400 12520
rect 37060 12880 38000 12900
rect 37060 12740 37080 12880
rect 37360 12740 37720 12880
rect 37980 12740 38000 12880
rect 37060 12660 38000 12740
rect 37060 12520 37080 12660
rect 37360 12520 37720 12660
rect 37980 12520 38000 12660
rect 37060 12500 38000 12520
rect 38660 12880 39600 12900
rect 38660 12740 38680 12880
rect 38960 12740 39320 12880
rect 39580 12740 39600 12880
rect 38660 12660 39600 12740
rect 38660 12520 38680 12660
rect 38960 12520 39320 12660
rect 39580 12520 39600 12660
rect 38660 12500 39600 12520
rect 40260 12880 41200 12900
rect 40260 12740 40280 12880
rect 40560 12740 40920 12880
rect 41180 12740 41200 12880
rect 40260 12660 41200 12740
rect 40260 12520 40280 12660
rect 40560 12520 40920 12660
rect 41180 12520 41200 12660
rect 40260 12500 41200 12520
rect 41860 12880 42800 12900
rect 41860 12740 41880 12880
rect 42160 12740 42520 12880
rect 42780 12740 42800 12880
rect 41860 12660 42800 12740
rect 41860 12520 41880 12660
rect 42160 12520 42520 12660
rect 42780 12520 42800 12660
rect 41860 12500 42800 12520
rect 43460 12880 44400 12900
rect 43460 12740 43480 12880
rect 43760 12740 44120 12880
rect 44380 12740 44400 12880
rect 43460 12660 44400 12740
rect 43460 12520 43480 12660
rect 43760 12520 44120 12660
rect 44380 12520 44400 12660
rect 43460 12500 44400 12520
rect 45060 12880 46000 12900
rect 45060 12740 45080 12880
rect 45360 12740 45720 12880
rect 45980 12740 46000 12880
rect 45060 12660 46000 12740
rect 45060 12520 45080 12660
rect 45360 12520 45720 12660
rect 45980 12520 46000 12660
rect 45060 12500 46000 12520
rect 46660 12880 47600 12900
rect 46660 12740 46680 12880
rect 46960 12740 47320 12880
rect 47580 12740 47600 12880
rect 46660 12660 47600 12740
rect 46660 12520 46680 12660
rect 46960 12520 47320 12660
rect 47580 12520 47600 12660
rect 46660 12500 47600 12520
rect 48260 12880 49200 12900
rect 48260 12740 48280 12880
rect 48560 12740 48920 12880
rect 49180 12740 49200 12880
rect 48260 12660 49200 12740
rect 48260 12520 48280 12660
rect 48560 12520 48920 12660
rect 49180 12520 49200 12660
rect 48260 12500 49200 12520
rect 49860 12880 50800 12900
rect 49860 12740 49880 12880
rect 50160 12740 50520 12880
rect 50780 12740 50800 12880
rect 49860 12660 50800 12740
rect 49860 12520 49880 12660
rect 50160 12520 50520 12660
rect 50780 12520 50800 12660
rect 49860 12500 50800 12520
rect 51460 12880 52400 12900
rect 51460 12740 51480 12880
rect 51760 12740 52120 12880
rect 52380 12740 52400 12880
rect 51460 12660 52400 12740
rect 51460 12520 51480 12660
rect 51760 12520 52120 12660
rect 52380 12520 52400 12660
rect 51460 12500 52400 12520
rect 53060 12880 54000 12900
rect 53060 12740 53080 12880
rect 53360 12740 53720 12880
rect 53980 12740 54000 12880
rect 53060 12660 54000 12740
rect 53060 12520 53080 12660
rect 53360 12520 53720 12660
rect 53980 12520 54000 12660
rect 53060 12500 54000 12520
rect 54660 12880 55600 12900
rect 54660 12740 54680 12880
rect 54960 12740 55320 12880
rect 55580 12740 55600 12880
rect 54660 12660 55600 12740
rect 54660 12520 54680 12660
rect 54960 12520 55320 12660
rect 55580 12520 55600 12660
rect 54660 12500 55600 12520
rect 56260 12880 57200 12900
rect 56260 12740 56280 12880
rect 56560 12740 56920 12880
rect 57180 12740 57200 12880
rect 56260 12660 57200 12740
rect 56260 12520 56280 12660
rect 56560 12520 56920 12660
rect 57180 12520 57200 12660
rect 56260 12500 57200 12520
rect 57860 12880 58800 12900
rect 57860 12740 57880 12880
rect 58160 12740 58520 12880
rect 58780 12740 58800 12880
rect 57860 12660 58800 12740
rect 57860 12520 57880 12660
rect 58160 12520 58520 12660
rect 58780 12520 58800 12660
rect 57860 12500 58800 12520
rect 59460 12880 60400 12900
rect 59460 12740 59480 12880
rect 59760 12740 60120 12880
rect 60380 12740 60400 12880
rect 59460 12660 60400 12740
rect 59460 12520 59480 12660
rect 59760 12520 60120 12660
rect 60380 12520 60400 12660
rect 59460 12500 60400 12520
rect 61060 12880 62000 12900
rect 61060 12740 61080 12880
rect 61360 12740 61720 12880
rect 61980 12740 62000 12880
rect 61060 12660 62000 12740
rect 61060 12520 61080 12660
rect 61360 12520 61720 12660
rect 61980 12520 62000 12660
rect 61060 12500 62000 12520
rect 62660 12880 63600 12900
rect 62660 12740 62680 12880
rect 62960 12740 63320 12880
rect 63580 12740 63600 12880
rect 62660 12660 63600 12740
rect 62660 12520 62680 12660
rect 62960 12520 63320 12660
rect 63580 12520 63600 12660
rect 62660 12500 63600 12520
rect 64260 12880 65200 12900
rect 64260 12740 64280 12880
rect 64560 12740 64920 12880
rect 65180 12740 65200 12880
rect 64260 12660 65200 12740
rect 64260 12520 64280 12660
rect 64560 12520 64920 12660
rect 65180 12520 65200 12660
rect 64260 12500 65200 12520
rect 65860 12880 66800 12900
rect 65860 12740 65880 12880
rect 66160 12740 66520 12880
rect 66780 12740 66800 12880
rect 65860 12660 66800 12740
rect 65860 12520 65880 12660
rect 66160 12520 66520 12660
rect 66780 12520 66800 12660
rect 65860 12500 66800 12520
rect 67460 12880 68400 12900
rect 67460 12740 67480 12880
rect 67760 12740 68120 12880
rect 68380 12740 68400 12880
rect 67460 12660 68400 12740
rect 67460 12520 67480 12660
rect 67760 12520 68120 12660
rect 68380 12520 68400 12660
rect 67460 12500 68400 12520
rect 69060 12880 70000 12900
rect 69060 12740 69080 12880
rect 69360 12740 69720 12880
rect 69980 12740 70000 12880
rect 69060 12660 70000 12740
rect 69060 12520 69080 12660
rect 69360 12520 69720 12660
rect 69980 12520 70000 12660
rect 69060 12500 70000 12520
rect 70660 12880 71600 12900
rect 70660 12740 70680 12880
rect 70960 12740 71320 12880
rect 71580 12740 71600 12880
rect 70660 12660 71600 12740
rect 70660 12520 70680 12660
rect 70960 12520 71320 12660
rect 71580 12520 71600 12660
rect 70660 12500 71600 12520
rect 72260 12880 73200 12900
rect 72260 12740 72280 12880
rect 72560 12740 72920 12880
rect 73180 12740 73200 12880
rect 72260 12660 73200 12740
rect 72260 12520 72280 12660
rect 72560 12520 72920 12660
rect 73180 12520 73200 12660
rect 72260 12500 73200 12520
rect 73860 12880 74800 12900
rect 73860 12740 73880 12880
rect 74160 12740 74520 12880
rect 74780 12740 74800 12880
rect 73860 12660 74800 12740
rect 73860 12520 73880 12660
rect 74160 12520 74520 12660
rect 74780 12520 74800 12660
rect 73860 12500 74800 12520
rect 75460 12880 76400 12900
rect 75460 12740 75480 12880
rect 75760 12740 76120 12880
rect 76380 12740 76400 12880
rect 75460 12660 76400 12740
rect 75460 12520 75480 12660
rect 75760 12520 76120 12660
rect 76380 12520 76400 12660
rect 75460 12500 76400 12520
rect 77060 12880 78000 12900
rect 77060 12740 77080 12880
rect 77360 12740 77720 12880
rect 77980 12740 78000 12880
rect 77060 12660 78000 12740
rect 77060 12520 77080 12660
rect 77360 12520 77720 12660
rect 77980 12520 78000 12660
rect 77060 12500 78000 12520
rect 78660 12880 79600 12900
rect 78660 12740 78680 12880
rect 78960 12740 79320 12880
rect 79580 12740 79600 12880
rect 78660 12660 79600 12740
rect 78660 12520 78680 12660
rect 78960 12520 79320 12660
rect 79580 12520 79600 12660
rect 78660 12500 79600 12520
rect 80260 12880 81200 12900
rect 80260 12740 80280 12880
rect 80560 12740 80920 12880
rect 81180 12740 81200 12880
rect 80260 12660 81200 12740
rect 80260 12520 80280 12660
rect 80560 12520 80920 12660
rect 81180 12520 81200 12660
rect 80260 12500 81200 12520
rect 81860 12880 82800 12900
rect 81860 12740 81880 12880
rect 82160 12740 82520 12880
rect 82780 12740 82800 12880
rect 81860 12660 82800 12740
rect 81860 12520 81880 12660
rect 82160 12520 82520 12660
rect 82780 12520 82800 12660
rect 81860 12500 82800 12520
rect 83460 12880 84400 12900
rect 83460 12740 83480 12880
rect 83760 12740 84120 12880
rect 84380 12740 84400 12880
rect 83460 12660 84400 12740
rect 83460 12520 83480 12660
rect 83760 12520 84120 12660
rect 84380 12520 84400 12660
rect 83460 12500 84400 12520
rect 85060 12880 86000 12900
rect 85060 12740 85080 12880
rect 85360 12740 85720 12880
rect 85980 12740 86000 12880
rect 85060 12660 86000 12740
rect 85060 12520 85080 12660
rect 85360 12520 85720 12660
rect 85980 12520 86000 12660
rect 85060 12500 86000 12520
rect 86660 12880 87600 12900
rect 86660 12740 86680 12880
rect 86960 12740 87320 12880
rect 87580 12740 87600 12880
rect 86660 12660 87600 12740
rect 86660 12520 86680 12660
rect 86960 12520 87320 12660
rect 87580 12520 87600 12660
rect 86660 12500 87600 12520
rect -33100 12380 -32680 12500
rect -33580 12220 -32680 12380
rect -33580 12080 -33540 12220
rect -33160 12180 -32680 12220
rect -33160 12080 -33100 12180
rect -33580 12040 -33100 12080
<< via3 >>
rect -33320 12740 -33040 12880
rect -32680 12740 -32420 12880
rect -33320 12520 -33040 12660
rect -32680 12520 -32420 12660
rect -31720 12740 -31440 12880
rect -31080 12740 -30820 12880
rect -31720 12520 -31440 12660
rect -31080 12520 -30820 12660
rect -30120 12740 -29840 12880
rect -29480 12740 -29220 12880
rect -30120 12520 -29840 12660
rect -29480 12520 -29220 12660
rect -28520 12740 -28240 12880
rect -27880 12740 -27620 12880
rect -28520 12520 -28240 12660
rect -27880 12520 -27620 12660
rect -26920 12740 -26640 12880
rect -26280 12740 -26020 12880
rect -26920 12520 -26640 12660
rect -26280 12520 -26020 12660
rect -25320 12740 -25040 12880
rect -24680 12740 -24420 12880
rect -25320 12520 -25040 12660
rect -24680 12520 -24420 12660
rect -23720 12740 -23440 12880
rect -23080 12740 -22820 12880
rect -23720 12520 -23440 12660
rect -23080 12520 -22820 12660
rect -22120 12740 -21840 12880
rect -21480 12740 -21220 12880
rect -22120 12520 -21840 12660
rect -21480 12520 -21220 12660
rect -20520 12740 -20240 12880
rect -19880 12740 -19620 12880
rect -20520 12520 -20240 12660
rect -19880 12520 -19620 12660
rect -18920 12740 -18640 12880
rect -18280 12740 -18020 12880
rect -18920 12520 -18640 12660
rect -18280 12520 -18020 12660
rect -17320 12740 -17040 12880
rect -16680 12740 -16420 12880
rect -17320 12520 -17040 12660
rect -16680 12520 -16420 12660
rect -15720 12740 -15440 12880
rect -15080 12740 -14820 12880
rect -15720 12520 -15440 12660
rect -15080 12520 -14820 12660
rect -14120 12740 -13840 12880
rect -13480 12740 -13220 12880
rect -14120 12520 -13840 12660
rect -13480 12520 -13220 12660
rect -12520 12740 -12240 12880
rect -11880 12740 -11620 12880
rect -12520 12520 -12240 12660
rect -11880 12520 -11620 12660
rect -10920 12740 -10640 12880
rect -10280 12740 -10020 12880
rect -10920 12520 -10640 12660
rect -10280 12520 -10020 12660
rect -9320 12740 -9040 12880
rect -8680 12740 -8420 12880
rect -9320 12520 -9040 12660
rect -8680 12520 -8420 12660
rect -7720 12740 -7440 12880
rect -7080 12740 -6820 12880
rect -7720 12520 -7440 12660
rect -7080 12520 -6820 12660
rect -6120 12740 -5840 12880
rect -5480 12740 -5220 12880
rect -6120 12520 -5840 12660
rect -5480 12520 -5220 12660
rect -4520 12740 -4240 12880
rect -3880 12740 -3620 12880
rect -4520 12520 -4240 12660
rect -3880 12520 -3620 12660
rect -2920 12740 -2640 12880
rect -2280 12740 -2020 12880
rect -2920 12520 -2640 12660
rect -2280 12520 -2020 12660
rect -1320 12740 -1040 12880
rect -680 12740 -420 12880
rect -1320 12520 -1040 12660
rect -680 12520 -420 12660
rect 280 12740 560 12880
rect 920 12740 1180 12880
rect 280 12520 560 12660
rect 920 12520 1180 12660
rect 1880 12740 2160 12880
rect 2520 12740 2780 12880
rect 1880 12520 2160 12660
rect 2520 12520 2780 12660
rect 3480 12740 3760 12880
rect 4120 12740 4380 12880
rect 3480 12520 3760 12660
rect 4120 12520 4380 12660
rect 5080 12740 5360 12880
rect 5720 12740 5980 12880
rect 5080 12520 5360 12660
rect 5720 12520 5980 12660
rect 6680 12740 6960 12880
rect 7320 12740 7580 12880
rect 6680 12520 6960 12660
rect 7320 12520 7580 12660
rect 8280 12740 8560 12880
rect 8920 12740 9180 12880
rect 8280 12520 8560 12660
rect 8920 12520 9180 12660
rect 9880 12740 10160 12880
rect 10520 12740 10780 12880
rect 9880 12520 10160 12660
rect 10520 12520 10780 12660
rect 11480 12740 11760 12880
rect 12120 12740 12380 12880
rect 11480 12520 11760 12660
rect 12120 12520 12380 12660
rect 13080 12740 13360 12880
rect 13720 12740 13980 12880
rect 13080 12520 13360 12660
rect 13720 12520 13980 12660
rect 14680 12740 14960 12880
rect 15320 12740 15580 12880
rect 14680 12520 14960 12660
rect 15320 12520 15580 12660
rect 16280 12740 16560 12880
rect 16920 12740 17180 12880
rect 16280 12520 16560 12660
rect 16920 12520 17180 12660
rect 17880 12740 18160 12880
rect 18520 12740 18780 12880
rect 17880 12520 18160 12660
rect 18520 12520 18780 12660
rect 19480 12740 19760 12880
rect 20120 12740 20380 12880
rect 19480 12520 19760 12660
rect 20120 12520 20380 12660
rect 21080 12740 21360 12880
rect 21720 12740 21980 12880
rect 21080 12520 21360 12660
rect 21720 12520 21980 12660
rect 22680 12740 22960 12880
rect 23320 12740 23580 12880
rect 22680 12520 22960 12660
rect 23320 12520 23580 12660
rect 24280 12740 24560 12880
rect 24920 12740 25180 12880
rect 24280 12520 24560 12660
rect 24920 12520 25180 12660
rect 25880 12740 26160 12880
rect 26520 12740 26780 12880
rect 25880 12520 26160 12660
rect 26520 12520 26780 12660
rect 27480 12740 27760 12880
rect 28120 12740 28380 12880
rect 27480 12520 27760 12660
rect 28120 12520 28380 12660
rect 29080 12740 29360 12880
rect 29720 12740 29980 12880
rect 29080 12520 29360 12660
rect 29720 12520 29980 12660
rect 30680 12740 30960 12880
rect 31320 12740 31580 12880
rect 30680 12520 30960 12660
rect 31320 12520 31580 12660
rect 32280 12740 32560 12880
rect 32920 12740 33180 12880
rect 32280 12520 32560 12660
rect 32920 12520 33180 12660
rect 33880 12740 34160 12880
rect 34520 12740 34780 12880
rect 33880 12520 34160 12660
rect 34520 12520 34780 12660
rect 35480 12740 35760 12880
rect 36120 12740 36380 12880
rect 35480 12520 35760 12660
rect 36120 12520 36380 12660
rect 37080 12740 37360 12880
rect 37720 12740 37980 12880
rect 37080 12520 37360 12660
rect 37720 12520 37980 12660
rect 38680 12740 38960 12880
rect 39320 12740 39580 12880
rect 38680 12520 38960 12660
rect 39320 12520 39580 12660
rect 40280 12740 40560 12880
rect 40920 12740 41180 12880
rect 40280 12520 40560 12660
rect 40920 12520 41180 12660
rect 41880 12740 42160 12880
rect 42520 12740 42780 12880
rect 41880 12520 42160 12660
rect 42520 12520 42780 12660
rect 43480 12740 43760 12880
rect 44120 12740 44380 12880
rect 43480 12520 43760 12660
rect 44120 12520 44380 12660
rect 45080 12740 45360 12880
rect 45720 12740 45980 12880
rect 45080 12520 45360 12660
rect 45720 12520 45980 12660
rect 46680 12740 46960 12880
rect 47320 12740 47580 12880
rect 46680 12520 46960 12660
rect 47320 12520 47580 12660
rect 48280 12740 48560 12880
rect 48920 12740 49180 12880
rect 48280 12520 48560 12660
rect 48920 12520 49180 12660
rect 49880 12740 50160 12880
rect 50520 12740 50780 12880
rect 49880 12520 50160 12660
rect 50520 12520 50780 12660
rect 51480 12740 51760 12880
rect 52120 12740 52380 12880
rect 51480 12520 51760 12660
rect 52120 12520 52380 12660
rect 53080 12740 53360 12880
rect 53720 12740 53980 12880
rect 53080 12520 53360 12660
rect 53720 12520 53980 12660
rect 54680 12740 54960 12880
rect 55320 12740 55580 12880
rect 54680 12520 54960 12660
rect 55320 12520 55580 12660
rect 56280 12740 56560 12880
rect 56920 12740 57180 12880
rect 56280 12520 56560 12660
rect 56920 12520 57180 12660
rect 57880 12740 58160 12880
rect 58520 12740 58780 12880
rect 57880 12520 58160 12660
rect 58520 12520 58780 12660
rect 59480 12740 59760 12880
rect 60120 12740 60380 12880
rect 59480 12520 59760 12660
rect 60120 12520 60380 12660
rect 61080 12740 61360 12880
rect 61720 12740 61980 12880
rect 61080 12520 61360 12660
rect 61720 12520 61980 12660
rect 62680 12740 62960 12880
rect 63320 12740 63580 12880
rect 62680 12520 62960 12660
rect 63320 12520 63580 12660
rect 64280 12740 64560 12880
rect 64920 12740 65180 12880
rect 64280 12520 64560 12660
rect 64920 12520 65180 12660
rect 65880 12740 66160 12880
rect 66520 12740 66780 12880
rect 65880 12520 66160 12660
rect 66520 12520 66780 12660
rect 67480 12740 67760 12880
rect 68120 12740 68380 12880
rect 67480 12520 67760 12660
rect 68120 12520 68380 12660
rect 69080 12740 69360 12880
rect 69720 12740 69980 12880
rect 69080 12520 69360 12660
rect 69720 12520 69980 12660
rect 70680 12740 70960 12880
rect 71320 12740 71580 12880
rect 70680 12520 70960 12660
rect 71320 12520 71580 12660
rect 72280 12740 72560 12880
rect 72920 12740 73180 12880
rect 72280 12520 72560 12660
rect 72920 12520 73180 12660
rect 73880 12740 74160 12880
rect 74520 12740 74780 12880
rect 73880 12520 74160 12660
rect 74520 12520 74780 12660
rect 75480 12740 75760 12880
rect 76120 12740 76380 12880
rect 75480 12520 75760 12660
rect 76120 12520 76380 12660
rect 77080 12740 77360 12880
rect 77720 12740 77980 12880
rect 77080 12520 77360 12660
rect 77720 12520 77980 12660
rect 78680 12740 78960 12880
rect 79320 12740 79580 12880
rect 78680 12520 78960 12660
rect 79320 12520 79580 12660
rect 80280 12740 80560 12880
rect 80920 12740 81180 12880
rect 80280 12520 80560 12660
rect 80920 12520 81180 12660
rect 81880 12740 82160 12880
rect 82520 12740 82780 12880
rect 81880 12520 82160 12660
rect 82520 12520 82780 12660
rect 83480 12740 83760 12880
rect 84120 12740 84380 12880
rect 83480 12520 83760 12660
rect 84120 12520 84380 12660
rect 85080 12740 85360 12880
rect 85720 12740 85980 12880
rect 85080 12520 85360 12660
rect 85720 12520 85980 12660
rect 86680 12740 86960 12880
rect 87320 12740 87580 12880
rect 86680 12520 86960 12660
rect 87320 12520 87580 12660
<< metal4 >>
rect -33820 12900 -33700 13000
rect -32220 12900 -32100 13000
rect -30620 12900 -30500 13000
rect -29020 12900 -28900 13000
rect -27420 12900 -27300 13000
rect -25820 12900 -25700 13000
rect -24220 12900 -24100 13000
rect -22620 12900 -22500 13000
rect -21020 12900 -20900 13000
rect -19420 12900 -19300 13000
rect -17820 12900 -17700 13000
rect -16220 12900 -16100 13000
rect -14620 12900 -14500 13000
rect -13020 12900 -12900 13000
rect -11420 12900 -11300 13000
rect -9820 12900 -9700 13000
rect -8220 12900 -8100 13000
rect -6620 12900 -6500 13000
rect -5020 12900 -4900 13000
rect -3420 12900 -3300 13000
rect -1820 12900 -1700 13000
rect -220 12900 -100 13000
rect 1380 12900 1500 13000
rect 2980 12900 3100 13000
rect 4580 12900 4700 13000
rect 6180 12900 6300 13000
rect 7780 12900 7900 13000
rect 9380 12900 9500 13000
rect 10980 12900 11100 13000
rect 12580 12900 12700 13000
rect 14180 12900 14300 13000
rect 15780 12900 15900 13000
rect 17380 12900 17500 13000
rect 18980 12900 19100 13000
rect 20580 12900 20700 13000
rect 22180 12900 22300 13000
rect 23780 12900 23900 13000
rect 25380 12900 25500 13000
rect 26980 12900 27100 13000
rect 28580 12900 28700 13000
rect 30180 12900 30300 13000
rect 31780 12900 31900 13000
rect 33380 12900 33500 13000
rect 34980 12900 35100 13000
rect 36580 12900 36700 13000
rect 38180 12900 38300 13000
rect 39780 12900 39900 13000
rect 41380 12900 41500 13000
rect 42980 12900 43100 13000
rect 44580 12900 44700 13000
rect 46180 12900 46300 13000
rect 47780 12900 47900 13000
rect 49380 12900 49500 13000
rect 50980 12900 51100 13000
rect 52580 12900 52700 13000
rect 54180 12900 54300 13000
rect 55780 12900 55900 13000
rect 57380 12900 57500 13000
rect 58980 12900 59100 13000
rect 60580 12900 60700 13000
rect 62180 12900 62300 13000
rect 63780 12900 63900 13000
rect 65380 12900 65500 13000
rect 66980 12900 67100 13000
rect 68580 12900 68700 13000
rect 70180 12900 70300 13000
rect 71780 12900 71900 13000
rect 73380 12900 73500 13000
rect 74980 12900 75100 13000
rect 76580 12900 76700 13000
rect 78180 12900 78300 13000
rect 79780 12900 79900 13000
rect 81380 12900 81500 13000
rect 82980 12900 83100 13000
rect 84580 12900 84700 13000
rect 86180 12900 86300 13000
rect -33820 12880 -33000 12900
rect -33820 12740 -33320 12880
rect -33040 12740 -33000 12880
rect -33820 12660 -33000 12740
rect -33820 12520 -33320 12660
rect -33040 12520 -33000 12660
rect -33820 12500 -33000 12520
rect -32700 12880 -31400 12900
rect -32700 12740 -32680 12880
rect -32420 12740 -31720 12880
rect -31440 12740 -31400 12880
rect -32700 12660 -31400 12740
rect -32700 12520 -32680 12660
rect -32420 12520 -31720 12660
rect -31440 12520 -31400 12660
rect -32700 12500 -31400 12520
rect -31100 12880 -29800 12900
rect -31100 12740 -31080 12880
rect -30820 12740 -30120 12880
rect -29840 12740 -29800 12880
rect -31100 12660 -29800 12740
rect -31100 12520 -31080 12660
rect -30820 12520 -30120 12660
rect -29840 12520 -29800 12660
rect -31100 12500 -29800 12520
rect -29500 12880 -28200 12900
rect -29500 12740 -29480 12880
rect -29220 12740 -28520 12880
rect -28240 12740 -28200 12880
rect -29500 12660 -28200 12740
rect -29500 12520 -29480 12660
rect -29220 12520 -28520 12660
rect -28240 12520 -28200 12660
rect -29500 12500 -28200 12520
rect -27900 12880 -26600 12900
rect -27900 12740 -27880 12880
rect -27620 12740 -26920 12880
rect -26640 12740 -26600 12880
rect -27900 12660 -26600 12740
rect -27900 12520 -27880 12660
rect -27620 12520 -26920 12660
rect -26640 12520 -26600 12660
rect -27900 12500 -26600 12520
rect -26300 12880 -25000 12900
rect -26300 12740 -26280 12880
rect -26020 12740 -25320 12880
rect -25040 12740 -25000 12880
rect -26300 12660 -25000 12740
rect -26300 12520 -26280 12660
rect -26020 12520 -25320 12660
rect -25040 12520 -25000 12660
rect -26300 12500 -25000 12520
rect -24700 12880 -23400 12900
rect -24700 12740 -24680 12880
rect -24420 12740 -23720 12880
rect -23440 12740 -23400 12880
rect -24700 12660 -23400 12740
rect -24700 12520 -24680 12660
rect -24420 12520 -23720 12660
rect -23440 12520 -23400 12660
rect -24700 12500 -23400 12520
rect -23100 12880 -21800 12900
rect -23100 12740 -23080 12880
rect -22820 12740 -22120 12880
rect -21840 12740 -21800 12880
rect -23100 12660 -21800 12740
rect -23100 12520 -23080 12660
rect -22820 12520 -22120 12660
rect -21840 12520 -21800 12660
rect -23100 12500 -21800 12520
rect -21500 12880 -20200 12900
rect -21500 12740 -21480 12880
rect -21220 12740 -20520 12880
rect -20240 12740 -20200 12880
rect -21500 12660 -20200 12740
rect -21500 12520 -21480 12660
rect -21220 12520 -20520 12660
rect -20240 12520 -20200 12660
rect -21500 12500 -20200 12520
rect -19900 12880 -18600 12900
rect -19900 12740 -19880 12880
rect -19620 12740 -18920 12880
rect -18640 12740 -18600 12880
rect -19900 12660 -18600 12740
rect -19900 12520 -19880 12660
rect -19620 12520 -18920 12660
rect -18640 12520 -18600 12660
rect -19900 12500 -18600 12520
rect -18300 12880 -17000 12900
rect -18300 12740 -18280 12880
rect -18020 12740 -17320 12880
rect -17040 12740 -17000 12880
rect -18300 12660 -17000 12740
rect -18300 12520 -18280 12660
rect -18020 12520 -17320 12660
rect -17040 12520 -17000 12660
rect -18300 12500 -17000 12520
rect -16700 12880 -15400 12900
rect -16700 12740 -16680 12880
rect -16420 12740 -15720 12880
rect -15440 12740 -15400 12880
rect -16700 12660 -15400 12740
rect -16700 12520 -16680 12660
rect -16420 12520 -15720 12660
rect -15440 12520 -15400 12660
rect -16700 12500 -15400 12520
rect -15100 12880 -13800 12900
rect -15100 12740 -15080 12880
rect -14820 12740 -14120 12880
rect -13840 12740 -13800 12880
rect -15100 12660 -13800 12740
rect -15100 12520 -15080 12660
rect -14820 12520 -14120 12660
rect -13840 12520 -13800 12660
rect -15100 12500 -13800 12520
rect -13500 12880 -12200 12900
rect -13500 12740 -13480 12880
rect -13220 12740 -12520 12880
rect -12240 12740 -12200 12880
rect -13500 12660 -12200 12740
rect -13500 12520 -13480 12660
rect -13220 12520 -12520 12660
rect -12240 12520 -12200 12660
rect -13500 12500 -12200 12520
rect -11900 12880 -10600 12900
rect -11900 12740 -11880 12880
rect -11620 12740 -10920 12880
rect -10640 12740 -10600 12880
rect -11900 12660 -10600 12740
rect -11900 12520 -11880 12660
rect -11620 12520 -10920 12660
rect -10640 12520 -10600 12660
rect -11900 12500 -10600 12520
rect -10300 12880 -9000 12900
rect -10300 12740 -10280 12880
rect -10020 12740 -9320 12880
rect -9040 12740 -9000 12880
rect -10300 12660 -9000 12740
rect -10300 12520 -10280 12660
rect -10020 12520 -9320 12660
rect -9040 12520 -9000 12660
rect -10300 12500 -9000 12520
rect -8700 12880 -7400 12900
rect -8700 12740 -8680 12880
rect -8420 12740 -7720 12880
rect -7440 12740 -7400 12880
rect -8700 12660 -7400 12740
rect -8700 12520 -8680 12660
rect -8420 12520 -7720 12660
rect -7440 12520 -7400 12660
rect -8700 12500 -7400 12520
rect -7100 12880 -5800 12900
rect -7100 12740 -7080 12880
rect -6820 12740 -6120 12880
rect -5840 12740 -5800 12880
rect -7100 12660 -5800 12740
rect -7100 12520 -7080 12660
rect -6820 12520 -6120 12660
rect -5840 12520 -5800 12660
rect -7100 12500 -5800 12520
rect -5500 12880 -4200 12900
rect -5500 12740 -5480 12880
rect -5220 12740 -4520 12880
rect -4240 12740 -4200 12880
rect -5500 12660 -4200 12740
rect -5500 12520 -5480 12660
rect -5220 12520 -4520 12660
rect -4240 12520 -4200 12660
rect -5500 12500 -4200 12520
rect -3900 12880 -2600 12900
rect -3900 12740 -3880 12880
rect -3620 12740 -2920 12880
rect -2640 12740 -2600 12880
rect -3900 12660 -2600 12740
rect -3900 12520 -3880 12660
rect -3620 12520 -2920 12660
rect -2640 12520 -2600 12660
rect -3900 12500 -2600 12520
rect -2300 12880 -1000 12900
rect -2300 12740 -2280 12880
rect -2020 12740 -1320 12880
rect -1040 12740 -1000 12880
rect -2300 12660 -1000 12740
rect -2300 12520 -2280 12660
rect -2020 12520 -1320 12660
rect -1040 12520 -1000 12660
rect -2300 12500 -1000 12520
rect -700 12880 600 12900
rect -700 12740 -680 12880
rect -420 12740 280 12880
rect 560 12740 600 12880
rect -700 12660 600 12740
rect -700 12520 -680 12660
rect -420 12520 280 12660
rect 560 12520 600 12660
rect -700 12500 600 12520
rect 900 12880 2200 12900
rect 900 12740 920 12880
rect 1180 12740 1880 12880
rect 2160 12740 2200 12880
rect 900 12660 2200 12740
rect 900 12520 920 12660
rect 1180 12520 1880 12660
rect 2160 12520 2200 12660
rect 900 12500 2200 12520
rect 2500 12880 3800 12900
rect 2500 12740 2520 12880
rect 2780 12740 3480 12880
rect 3760 12740 3800 12880
rect 2500 12660 3800 12740
rect 2500 12520 2520 12660
rect 2780 12520 3480 12660
rect 3760 12520 3800 12660
rect 2500 12500 3800 12520
rect 4100 12880 5400 12900
rect 4100 12740 4120 12880
rect 4380 12740 5080 12880
rect 5360 12740 5400 12880
rect 4100 12660 5400 12740
rect 4100 12520 4120 12660
rect 4380 12520 5080 12660
rect 5360 12520 5400 12660
rect 4100 12500 5400 12520
rect 5700 12880 7000 12900
rect 5700 12740 5720 12880
rect 5980 12740 6680 12880
rect 6960 12740 7000 12880
rect 5700 12660 7000 12740
rect 5700 12520 5720 12660
rect 5980 12520 6680 12660
rect 6960 12520 7000 12660
rect 5700 12500 7000 12520
rect 7300 12880 8600 12900
rect 7300 12740 7320 12880
rect 7580 12740 8280 12880
rect 8560 12740 8600 12880
rect 7300 12660 8600 12740
rect 7300 12520 7320 12660
rect 7580 12520 8280 12660
rect 8560 12520 8600 12660
rect 7300 12500 8600 12520
rect 8900 12880 10200 12900
rect 8900 12740 8920 12880
rect 9180 12740 9880 12880
rect 10160 12740 10200 12880
rect 8900 12660 10200 12740
rect 8900 12520 8920 12660
rect 9180 12520 9880 12660
rect 10160 12520 10200 12660
rect 8900 12500 10200 12520
rect 10500 12880 11800 12900
rect 10500 12740 10520 12880
rect 10780 12740 11480 12880
rect 11760 12740 11800 12880
rect 10500 12660 11800 12740
rect 10500 12520 10520 12660
rect 10780 12520 11480 12660
rect 11760 12520 11800 12660
rect 10500 12500 11800 12520
rect 12100 12880 13400 12900
rect 12100 12740 12120 12880
rect 12380 12740 13080 12880
rect 13360 12740 13400 12880
rect 12100 12660 13400 12740
rect 12100 12520 12120 12660
rect 12380 12520 13080 12660
rect 13360 12520 13400 12660
rect 12100 12500 13400 12520
rect 13700 12880 15000 12900
rect 13700 12740 13720 12880
rect 13980 12740 14680 12880
rect 14960 12740 15000 12880
rect 13700 12660 15000 12740
rect 13700 12520 13720 12660
rect 13980 12520 14680 12660
rect 14960 12520 15000 12660
rect 13700 12500 15000 12520
rect 15300 12880 16600 12900
rect 15300 12740 15320 12880
rect 15580 12740 16280 12880
rect 16560 12740 16600 12880
rect 15300 12660 16600 12740
rect 15300 12520 15320 12660
rect 15580 12520 16280 12660
rect 16560 12520 16600 12660
rect 15300 12500 16600 12520
rect 16900 12880 18200 12900
rect 16900 12740 16920 12880
rect 17180 12740 17880 12880
rect 18160 12740 18200 12880
rect 16900 12660 18200 12740
rect 16900 12520 16920 12660
rect 17180 12520 17880 12660
rect 18160 12520 18200 12660
rect 16900 12500 18200 12520
rect 18500 12880 19800 12900
rect 18500 12740 18520 12880
rect 18780 12740 19480 12880
rect 19760 12740 19800 12880
rect 18500 12660 19800 12740
rect 18500 12520 18520 12660
rect 18780 12520 19480 12660
rect 19760 12520 19800 12660
rect 18500 12500 19800 12520
rect 20100 12880 21400 12900
rect 20100 12740 20120 12880
rect 20380 12740 21080 12880
rect 21360 12740 21400 12880
rect 20100 12660 21400 12740
rect 20100 12520 20120 12660
rect 20380 12520 21080 12660
rect 21360 12520 21400 12660
rect 20100 12500 21400 12520
rect 21700 12880 23000 12900
rect 21700 12740 21720 12880
rect 21980 12740 22680 12880
rect 22960 12740 23000 12880
rect 21700 12660 23000 12740
rect 21700 12520 21720 12660
rect 21980 12520 22680 12660
rect 22960 12520 23000 12660
rect 21700 12500 23000 12520
rect 23300 12880 24600 12900
rect 23300 12740 23320 12880
rect 23580 12740 24280 12880
rect 24560 12740 24600 12880
rect 23300 12660 24600 12740
rect 23300 12520 23320 12660
rect 23580 12520 24280 12660
rect 24560 12520 24600 12660
rect 23300 12500 24600 12520
rect 24900 12880 26200 12900
rect 24900 12740 24920 12880
rect 25180 12740 25880 12880
rect 26160 12740 26200 12880
rect 24900 12660 26200 12740
rect 24900 12520 24920 12660
rect 25180 12520 25880 12660
rect 26160 12520 26200 12660
rect 24900 12500 26200 12520
rect 26500 12880 27800 12900
rect 26500 12740 26520 12880
rect 26780 12740 27480 12880
rect 27760 12740 27800 12880
rect 26500 12660 27800 12740
rect 26500 12520 26520 12660
rect 26780 12520 27480 12660
rect 27760 12520 27800 12660
rect 26500 12500 27800 12520
rect 28100 12880 29400 12900
rect 28100 12740 28120 12880
rect 28380 12740 29080 12880
rect 29360 12740 29400 12880
rect 28100 12660 29400 12740
rect 28100 12520 28120 12660
rect 28380 12520 29080 12660
rect 29360 12520 29400 12660
rect 28100 12500 29400 12520
rect 29700 12880 31000 12900
rect 29700 12740 29720 12880
rect 29980 12740 30680 12880
rect 30960 12740 31000 12880
rect 29700 12660 31000 12740
rect 29700 12520 29720 12660
rect 29980 12520 30680 12660
rect 30960 12520 31000 12660
rect 29700 12500 31000 12520
rect 31300 12880 32600 12900
rect 31300 12740 31320 12880
rect 31580 12740 32280 12880
rect 32560 12740 32600 12880
rect 31300 12660 32600 12740
rect 31300 12520 31320 12660
rect 31580 12520 32280 12660
rect 32560 12520 32600 12660
rect 31300 12500 32600 12520
rect 32900 12880 34200 12900
rect 32900 12740 32920 12880
rect 33180 12740 33880 12880
rect 34160 12740 34200 12880
rect 32900 12660 34200 12740
rect 32900 12520 32920 12660
rect 33180 12520 33880 12660
rect 34160 12520 34200 12660
rect 32900 12500 34200 12520
rect 34500 12880 35800 12900
rect 34500 12740 34520 12880
rect 34780 12740 35480 12880
rect 35760 12740 35800 12880
rect 34500 12660 35800 12740
rect 34500 12520 34520 12660
rect 34780 12520 35480 12660
rect 35760 12520 35800 12660
rect 34500 12500 35800 12520
rect 36100 12880 37400 12900
rect 36100 12740 36120 12880
rect 36380 12740 37080 12880
rect 37360 12740 37400 12880
rect 36100 12660 37400 12740
rect 36100 12520 36120 12660
rect 36380 12520 37080 12660
rect 37360 12520 37400 12660
rect 36100 12500 37400 12520
rect 37700 12880 39000 12900
rect 37700 12740 37720 12880
rect 37980 12740 38680 12880
rect 38960 12740 39000 12880
rect 37700 12660 39000 12740
rect 37700 12520 37720 12660
rect 37980 12520 38680 12660
rect 38960 12520 39000 12660
rect 37700 12500 39000 12520
rect 39300 12880 40600 12900
rect 39300 12740 39320 12880
rect 39580 12740 40280 12880
rect 40560 12740 40600 12880
rect 39300 12660 40600 12740
rect 39300 12520 39320 12660
rect 39580 12520 40280 12660
rect 40560 12520 40600 12660
rect 39300 12500 40600 12520
rect 40900 12880 42200 12900
rect 40900 12740 40920 12880
rect 41180 12740 41880 12880
rect 42160 12740 42200 12880
rect 40900 12660 42200 12740
rect 40900 12520 40920 12660
rect 41180 12520 41880 12660
rect 42160 12520 42200 12660
rect 40900 12500 42200 12520
rect 42500 12880 43800 12900
rect 42500 12740 42520 12880
rect 42780 12740 43480 12880
rect 43760 12740 43800 12880
rect 42500 12660 43800 12740
rect 42500 12520 42520 12660
rect 42780 12520 43480 12660
rect 43760 12520 43800 12660
rect 42500 12500 43800 12520
rect 44100 12880 45400 12900
rect 44100 12740 44120 12880
rect 44380 12740 45080 12880
rect 45360 12740 45400 12880
rect 44100 12660 45400 12740
rect 44100 12520 44120 12660
rect 44380 12520 45080 12660
rect 45360 12520 45400 12660
rect 44100 12500 45400 12520
rect 45700 12880 47000 12900
rect 45700 12740 45720 12880
rect 45980 12740 46680 12880
rect 46960 12740 47000 12880
rect 45700 12660 47000 12740
rect 45700 12520 45720 12660
rect 45980 12520 46680 12660
rect 46960 12520 47000 12660
rect 45700 12500 47000 12520
rect 47300 12880 48600 12900
rect 47300 12740 47320 12880
rect 47580 12740 48280 12880
rect 48560 12740 48600 12880
rect 47300 12660 48600 12740
rect 47300 12520 47320 12660
rect 47580 12520 48280 12660
rect 48560 12520 48600 12660
rect 47300 12500 48600 12520
rect 48900 12880 50200 12900
rect 48900 12740 48920 12880
rect 49180 12740 49880 12880
rect 50160 12740 50200 12880
rect 48900 12660 50200 12740
rect 48900 12520 48920 12660
rect 49180 12520 49880 12660
rect 50160 12520 50200 12660
rect 48900 12500 50200 12520
rect 50500 12880 51800 12900
rect 50500 12740 50520 12880
rect 50780 12740 51480 12880
rect 51760 12740 51800 12880
rect 50500 12660 51800 12740
rect 50500 12520 50520 12660
rect 50780 12520 51480 12660
rect 51760 12520 51800 12660
rect 50500 12500 51800 12520
rect 52100 12880 53400 12900
rect 52100 12740 52120 12880
rect 52380 12740 53080 12880
rect 53360 12740 53400 12880
rect 52100 12660 53400 12740
rect 52100 12520 52120 12660
rect 52380 12520 53080 12660
rect 53360 12520 53400 12660
rect 52100 12500 53400 12520
rect 53700 12880 55000 12900
rect 53700 12740 53720 12880
rect 53980 12740 54680 12880
rect 54960 12740 55000 12880
rect 53700 12660 55000 12740
rect 53700 12520 53720 12660
rect 53980 12520 54680 12660
rect 54960 12520 55000 12660
rect 53700 12500 55000 12520
rect 55300 12880 56600 12900
rect 55300 12740 55320 12880
rect 55580 12740 56280 12880
rect 56560 12740 56600 12880
rect 55300 12660 56600 12740
rect 55300 12520 55320 12660
rect 55580 12520 56280 12660
rect 56560 12520 56600 12660
rect 55300 12500 56600 12520
rect 56900 12880 58200 12900
rect 56900 12740 56920 12880
rect 57180 12740 57880 12880
rect 58160 12740 58200 12880
rect 56900 12660 58200 12740
rect 56900 12520 56920 12660
rect 57180 12520 57880 12660
rect 58160 12520 58200 12660
rect 56900 12500 58200 12520
rect 58500 12880 59800 12900
rect 58500 12740 58520 12880
rect 58780 12740 59480 12880
rect 59760 12740 59800 12880
rect 58500 12660 59800 12740
rect 58500 12520 58520 12660
rect 58780 12520 59480 12660
rect 59760 12520 59800 12660
rect 58500 12500 59800 12520
rect 60100 12880 61400 12900
rect 60100 12740 60120 12880
rect 60380 12740 61080 12880
rect 61360 12740 61400 12880
rect 60100 12660 61400 12740
rect 60100 12520 60120 12660
rect 60380 12520 61080 12660
rect 61360 12520 61400 12660
rect 60100 12500 61400 12520
rect 61700 12880 63000 12900
rect 61700 12740 61720 12880
rect 61980 12740 62680 12880
rect 62960 12740 63000 12880
rect 61700 12660 63000 12740
rect 61700 12520 61720 12660
rect 61980 12520 62680 12660
rect 62960 12520 63000 12660
rect 61700 12500 63000 12520
rect 63300 12880 64600 12900
rect 63300 12740 63320 12880
rect 63580 12740 64280 12880
rect 64560 12740 64600 12880
rect 63300 12660 64600 12740
rect 63300 12520 63320 12660
rect 63580 12520 64280 12660
rect 64560 12520 64600 12660
rect 63300 12500 64600 12520
rect 64900 12880 66200 12900
rect 64900 12740 64920 12880
rect 65180 12740 65880 12880
rect 66160 12740 66200 12880
rect 64900 12660 66200 12740
rect 64900 12520 64920 12660
rect 65180 12520 65880 12660
rect 66160 12520 66200 12660
rect 64900 12500 66200 12520
rect 66500 12880 67800 12900
rect 66500 12740 66520 12880
rect 66780 12740 67480 12880
rect 67760 12740 67800 12880
rect 66500 12660 67800 12740
rect 66500 12520 66520 12660
rect 66780 12520 67480 12660
rect 67760 12520 67800 12660
rect 66500 12500 67800 12520
rect 68100 12880 69400 12900
rect 68100 12740 68120 12880
rect 68380 12740 69080 12880
rect 69360 12740 69400 12880
rect 68100 12660 69400 12740
rect 68100 12520 68120 12660
rect 68380 12520 69080 12660
rect 69360 12520 69400 12660
rect 68100 12500 69400 12520
rect 69700 12880 71000 12900
rect 69700 12740 69720 12880
rect 69980 12740 70680 12880
rect 70960 12740 71000 12880
rect 69700 12660 71000 12740
rect 69700 12520 69720 12660
rect 69980 12520 70680 12660
rect 70960 12520 71000 12660
rect 69700 12500 71000 12520
rect 71300 12880 72600 12900
rect 71300 12740 71320 12880
rect 71580 12740 72280 12880
rect 72560 12740 72600 12880
rect 71300 12660 72600 12740
rect 71300 12520 71320 12660
rect 71580 12520 72280 12660
rect 72560 12520 72600 12660
rect 71300 12500 72600 12520
rect 72900 12880 74200 12900
rect 72900 12740 72920 12880
rect 73180 12740 73880 12880
rect 74160 12740 74200 12880
rect 72900 12660 74200 12740
rect 72900 12520 72920 12660
rect 73180 12520 73880 12660
rect 74160 12520 74200 12660
rect 72900 12500 74200 12520
rect 74500 12880 75800 12900
rect 74500 12740 74520 12880
rect 74780 12740 75480 12880
rect 75760 12740 75800 12880
rect 74500 12660 75800 12740
rect 74500 12520 74520 12660
rect 74780 12520 75480 12660
rect 75760 12520 75800 12660
rect 74500 12500 75800 12520
rect 76100 12880 77400 12900
rect 76100 12740 76120 12880
rect 76380 12740 77080 12880
rect 77360 12740 77400 12880
rect 76100 12660 77400 12740
rect 76100 12520 76120 12660
rect 76380 12520 77080 12660
rect 77360 12520 77400 12660
rect 76100 12500 77400 12520
rect 77700 12880 79000 12900
rect 77700 12740 77720 12880
rect 77980 12740 78680 12880
rect 78960 12740 79000 12880
rect 77700 12660 79000 12740
rect 77700 12520 77720 12660
rect 77980 12520 78680 12660
rect 78960 12520 79000 12660
rect 77700 12500 79000 12520
rect 79300 12880 80600 12900
rect 79300 12740 79320 12880
rect 79580 12740 80280 12880
rect 80560 12740 80600 12880
rect 79300 12660 80600 12740
rect 79300 12520 79320 12660
rect 79580 12520 80280 12660
rect 80560 12520 80600 12660
rect 79300 12500 80600 12520
rect 80900 12880 82200 12900
rect 80900 12740 80920 12880
rect 81180 12740 81880 12880
rect 82160 12740 82200 12880
rect 80900 12660 82200 12740
rect 80900 12520 80920 12660
rect 81180 12520 81880 12660
rect 82160 12520 82200 12660
rect 80900 12500 82200 12520
rect 82500 12880 83800 12900
rect 82500 12740 82520 12880
rect 82780 12740 83480 12880
rect 83760 12740 83800 12880
rect 82500 12660 83800 12740
rect 82500 12520 82520 12660
rect 82780 12520 83480 12660
rect 83760 12520 83800 12660
rect 82500 12500 83800 12520
rect 84100 12880 85400 12900
rect 84100 12740 84120 12880
rect 84380 12740 85080 12880
rect 85360 12740 85400 12880
rect 84100 12660 85400 12740
rect 84100 12520 84120 12660
rect 84380 12520 85080 12660
rect 85360 12520 85400 12660
rect 84100 12500 85400 12520
rect 85700 12880 87000 12900
rect 85700 12740 85720 12880
rect 85980 12740 86680 12880
rect 86960 12740 87000 12880
rect 85700 12660 87000 12740
rect 85700 12520 85720 12660
rect 85980 12520 86680 12660
rect 86960 12520 87000 12660
rect 85700 12500 87000 12520
rect 87300 12880 87780 12900
rect 87300 12740 87320 12880
rect 87580 12740 87780 12880
rect 87300 12660 87780 12740
rect 87300 12520 87320 12660
rect 87580 12520 87780 12660
rect 87300 12500 87780 12520
use cap1  cap1_0
timestamp 1667663783
transform 1 0 73800 0 1 13000
box 0 0 1300 1200
use cap1  cap1_4
timestamp 1667663783
transform 1 0 86600 0 1 13000
box 0 0 1300 1200
use cap1  cap1_5
timestamp 1667663783
transform 1 0 85000 0 1 13000
box 0 0 1300 1200
use cap2  cap2_0
timestamp 1667663783
transform 1 0 70600 0 1 13000
box 0 0 2900 1200
use cap2  cap2_3
timestamp 1667663783
transform 1 0 81800 0 1 13000
box 0 0 2900 1200
use cap4  cap4_0
timestamp 1667663783
transform 1 0 64200 0 1 13000
box 0 0 6100 1200
use cap4  cap4_1
timestamp 1667663783
transform 1 0 75400 0 1 13000
box 0 0 6100 1200
use cap8  cap8_0
timestamp 1667684479
transform 1 0 51400 0 1 13000
box 0 0 1300 12400
use cap8  cap8_1
timestamp 1667684479
transform 1 0 62600 0 1 13000
box 0 0 1300 12400
use cap16  cap16_0
timestamp 1667684462
transform 1 0 48200 0 1 13000
box 0 0 2900 12400
use cap16  cap16_1
timestamp 1667684462
transform 1 0 59400 0 1 13000
box 0 0 2900 12400
use cap32  cap32_0
timestamp 1667684412
transform 1 0 41800 0 1 13000
box 0 0 6100 12400
use cap32  cap32_1
timestamp 1667684412
transform 1 0 53000 0 1 13000
box 0 0 6100 12400
use cap64  cap64_0
timestamp 1667684360
transform 1 0 29000 0 1 13000
box 0 0 12500 12400
use cap64  cap64_1
timestamp 1667684360
transform 1 0 -9400 0 1 13000
box 0 0 12500 12400
use cap128  cap128_0
timestamp 1667663783
transform 1 0 -35000 0 1 13000
box 0 0 25300 12400
use cap128  cap128_1
timestamp 1667663783
transform 1 0 3400 0 1 13000
box 0 0 25300 12400
use sky130_fd_pr__nfet_01v8_HA267C  sky130_fd_pr__nfet_01v8_HA267C_0
timestamp 1667526910
transform 1 0 -33342 0 1 11057
box -258 -1057 258 1057
<< end >>
