magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -386 289772 386 289800
rect -386 285538 302 289772
rect 366 285538 386 289772
rect -386 285510 386 285538
rect -386 285242 386 285270
rect -386 281008 302 285242
rect 366 281008 386 285242
rect -386 280980 386 281008
rect -386 280712 386 280740
rect -386 276478 302 280712
rect 366 276478 386 280712
rect -386 276450 386 276478
rect -386 276182 386 276210
rect -386 271948 302 276182
rect 366 271948 386 276182
rect -386 271920 386 271948
rect -386 271652 386 271680
rect -386 267418 302 271652
rect 366 267418 386 271652
rect -386 267390 386 267418
rect -386 267122 386 267150
rect -386 262888 302 267122
rect 366 262888 386 267122
rect -386 262860 386 262888
rect -386 262592 386 262620
rect -386 258358 302 262592
rect 366 258358 386 262592
rect -386 258330 386 258358
rect -386 258062 386 258090
rect -386 253828 302 258062
rect 366 253828 386 258062
rect -386 253800 386 253828
rect -386 253532 386 253560
rect -386 249298 302 253532
rect 366 249298 386 253532
rect -386 249270 386 249298
rect -386 249002 386 249030
rect -386 244768 302 249002
rect 366 244768 386 249002
rect -386 244740 386 244768
rect -386 244472 386 244500
rect -386 240238 302 244472
rect 366 240238 386 244472
rect -386 240210 386 240238
rect -386 239942 386 239970
rect -386 235708 302 239942
rect 366 235708 386 239942
rect -386 235680 386 235708
rect -386 235412 386 235440
rect -386 231178 302 235412
rect 366 231178 386 235412
rect -386 231150 386 231178
rect -386 230882 386 230910
rect -386 226648 302 230882
rect 366 226648 386 230882
rect -386 226620 386 226648
rect -386 226352 386 226380
rect -386 222118 302 226352
rect 366 222118 386 226352
rect -386 222090 386 222118
rect -386 221822 386 221850
rect -386 217588 302 221822
rect 366 217588 386 221822
rect -386 217560 386 217588
rect -386 217292 386 217320
rect -386 213058 302 217292
rect 366 213058 386 217292
rect -386 213030 386 213058
rect -386 212762 386 212790
rect -386 208528 302 212762
rect 366 208528 386 212762
rect -386 208500 386 208528
rect -386 208232 386 208260
rect -386 203998 302 208232
rect 366 203998 386 208232
rect -386 203970 386 203998
rect -386 203702 386 203730
rect -386 199468 302 203702
rect 366 199468 386 203702
rect -386 199440 386 199468
rect -386 199172 386 199200
rect -386 194938 302 199172
rect 366 194938 386 199172
rect -386 194910 386 194938
rect -386 194642 386 194670
rect -386 190408 302 194642
rect 366 190408 386 194642
rect -386 190380 386 190408
rect -386 190112 386 190140
rect -386 185878 302 190112
rect 366 185878 386 190112
rect -386 185850 386 185878
rect -386 185582 386 185610
rect -386 181348 302 185582
rect 366 181348 386 185582
rect -386 181320 386 181348
rect -386 181052 386 181080
rect -386 176818 302 181052
rect 366 176818 386 181052
rect -386 176790 386 176818
rect -386 176522 386 176550
rect -386 172288 302 176522
rect 366 172288 386 176522
rect -386 172260 386 172288
rect -386 171992 386 172020
rect -386 167758 302 171992
rect 366 167758 386 171992
rect -386 167730 386 167758
rect -386 167462 386 167490
rect -386 163228 302 167462
rect 366 163228 386 167462
rect -386 163200 386 163228
rect -386 162932 386 162960
rect -386 158698 302 162932
rect 366 158698 386 162932
rect -386 158670 386 158698
rect -386 158402 386 158430
rect -386 154168 302 158402
rect 366 154168 386 158402
rect -386 154140 386 154168
rect -386 153872 386 153900
rect -386 149638 302 153872
rect 366 149638 386 153872
rect -386 149610 386 149638
rect -386 149342 386 149370
rect -386 145108 302 149342
rect 366 145108 386 149342
rect -386 145080 386 145108
rect -386 144812 386 144840
rect -386 140578 302 144812
rect 366 140578 386 144812
rect -386 140550 386 140578
rect -386 140282 386 140310
rect -386 136048 302 140282
rect 366 136048 386 140282
rect -386 136020 386 136048
rect -386 135752 386 135780
rect -386 131518 302 135752
rect 366 131518 386 135752
rect -386 131490 386 131518
rect -386 131222 386 131250
rect -386 126988 302 131222
rect 366 126988 386 131222
rect -386 126960 386 126988
rect -386 126692 386 126720
rect -386 122458 302 126692
rect 366 122458 386 126692
rect -386 122430 386 122458
rect -386 122162 386 122190
rect -386 117928 302 122162
rect 366 117928 386 122162
rect -386 117900 386 117928
rect -386 117632 386 117660
rect -386 113398 302 117632
rect 366 113398 386 117632
rect -386 113370 386 113398
rect -386 113102 386 113130
rect -386 108868 302 113102
rect 366 108868 386 113102
rect -386 108840 386 108868
rect -386 108572 386 108600
rect -386 104338 302 108572
rect 366 104338 386 108572
rect -386 104310 386 104338
rect -386 104042 386 104070
rect -386 99808 302 104042
rect 366 99808 386 104042
rect -386 99780 386 99808
rect -386 99512 386 99540
rect -386 95278 302 99512
rect 366 95278 386 99512
rect -386 95250 386 95278
rect -386 94982 386 95010
rect -386 90748 302 94982
rect 366 90748 386 94982
rect -386 90720 386 90748
rect -386 90452 386 90480
rect -386 86218 302 90452
rect 366 86218 386 90452
rect -386 86190 386 86218
rect -386 85922 386 85950
rect -386 81688 302 85922
rect 366 81688 386 85922
rect -386 81660 386 81688
rect -386 81392 386 81420
rect -386 77158 302 81392
rect 366 77158 386 81392
rect -386 77130 386 77158
rect -386 76862 386 76890
rect -386 72628 302 76862
rect 366 72628 386 76862
rect -386 72600 386 72628
rect -386 72332 386 72360
rect -386 68098 302 72332
rect 366 68098 386 72332
rect -386 68070 386 68098
rect -386 67802 386 67830
rect -386 63568 302 67802
rect 366 63568 386 67802
rect -386 63540 386 63568
rect -386 63272 386 63300
rect -386 59038 302 63272
rect 366 59038 386 63272
rect -386 59010 386 59038
rect -386 58742 386 58770
rect -386 54508 302 58742
rect 366 54508 386 58742
rect -386 54480 386 54508
rect -386 54212 386 54240
rect -386 49978 302 54212
rect 366 49978 386 54212
rect -386 49950 386 49978
rect -386 49682 386 49710
rect -386 45448 302 49682
rect 366 45448 386 49682
rect -386 45420 386 45448
rect -386 45152 386 45180
rect -386 40918 302 45152
rect 366 40918 386 45152
rect -386 40890 386 40918
rect -386 40622 386 40650
rect -386 36388 302 40622
rect 366 36388 386 40622
rect -386 36360 386 36388
rect -386 36092 386 36120
rect -386 31858 302 36092
rect 366 31858 386 36092
rect -386 31830 386 31858
rect -386 31562 386 31590
rect -386 27328 302 31562
rect 366 27328 386 31562
rect -386 27300 386 27328
rect -386 27032 386 27060
rect -386 22798 302 27032
rect 366 22798 386 27032
rect -386 22770 386 22798
rect -386 22502 386 22530
rect -386 18268 302 22502
rect 366 18268 386 22502
rect -386 18240 386 18268
rect -386 17972 386 18000
rect -386 13738 302 17972
rect 366 13738 386 17972
rect -386 13710 386 13738
rect -386 13442 386 13470
rect -386 9208 302 13442
rect 366 9208 386 13442
rect -386 9180 386 9208
rect -386 8912 386 8940
rect -386 4678 302 8912
rect 366 4678 386 8912
rect -386 4650 386 4678
rect -386 4382 386 4410
rect -386 148 302 4382
rect 366 148 386 4382
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -4382 302 -148
rect 366 -4382 386 -148
rect -386 -4410 386 -4382
rect -386 -4678 386 -4650
rect -386 -8912 302 -4678
rect 366 -8912 386 -4678
rect -386 -8940 386 -8912
rect -386 -9208 386 -9180
rect -386 -13442 302 -9208
rect 366 -13442 386 -9208
rect -386 -13470 386 -13442
rect -386 -13738 386 -13710
rect -386 -17972 302 -13738
rect 366 -17972 386 -13738
rect -386 -18000 386 -17972
rect -386 -18268 386 -18240
rect -386 -22502 302 -18268
rect 366 -22502 386 -18268
rect -386 -22530 386 -22502
rect -386 -22798 386 -22770
rect -386 -27032 302 -22798
rect 366 -27032 386 -22798
rect -386 -27060 386 -27032
rect -386 -27328 386 -27300
rect -386 -31562 302 -27328
rect 366 -31562 386 -27328
rect -386 -31590 386 -31562
rect -386 -31858 386 -31830
rect -386 -36092 302 -31858
rect 366 -36092 386 -31858
rect -386 -36120 386 -36092
rect -386 -36388 386 -36360
rect -386 -40622 302 -36388
rect 366 -40622 386 -36388
rect -386 -40650 386 -40622
rect -386 -40918 386 -40890
rect -386 -45152 302 -40918
rect 366 -45152 386 -40918
rect -386 -45180 386 -45152
rect -386 -45448 386 -45420
rect -386 -49682 302 -45448
rect 366 -49682 386 -45448
rect -386 -49710 386 -49682
rect -386 -49978 386 -49950
rect -386 -54212 302 -49978
rect 366 -54212 386 -49978
rect -386 -54240 386 -54212
rect -386 -54508 386 -54480
rect -386 -58742 302 -54508
rect 366 -58742 386 -54508
rect -386 -58770 386 -58742
rect -386 -59038 386 -59010
rect -386 -63272 302 -59038
rect 366 -63272 386 -59038
rect -386 -63300 386 -63272
rect -386 -63568 386 -63540
rect -386 -67802 302 -63568
rect 366 -67802 386 -63568
rect -386 -67830 386 -67802
rect -386 -68098 386 -68070
rect -386 -72332 302 -68098
rect 366 -72332 386 -68098
rect -386 -72360 386 -72332
rect -386 -72628 386 -72600
rect -386 -76862 302 -72628
rect 366 -76862 386 -72628
rect -386 -76890 386 -76862
rect -386 -77158 386 -77130
rect -386 -81392 302 -77158
rect 366 -81392 386 -77158
rect -386 -81420 386 -81392
rect -386 -81688 386 -81660
rect -386 -85922 302 -81688
rect 366 -85922 386 -81688
rect -386 -85950 386 -85922
rect -386 -86218 386 -86190
rect -386 -90452 302 -86218
rect 366 -90452 386 -86218
rect -386 -90480 386 -90452
rect -386 -90748 386 -90720
rect -386 -94982 302 -90748
rect 366 -94982 386 -90748
rect -386 -95010 386 -94982
rect -386 -95278 386 -95250
rect -386 -99512 302 -95278
rect 366 -99512 386 -95278
rect -386 -99540 386 -99512
rect -386 -99808 386 -99780
rect -386 -104042 302 -99808
rect 366 -104042 386 -99808
rect -386 -104070 386 -104042
rect -386 -104338 386 -104310
rect -386 -108572 302 -104338
rect 366 -108572 386 -104338
rect -386 -108600 386 -108572
rect -386 -108868 386 -108840
rect -386 -113102 302 -108868
rect 366 -113102 386 -108868
rect -386 -113130 386 -113102
rect -386 -113398 386 -113370
rect -386 -117632 302 -113398
rect 366 -117632 386 -113398
rect -386 -117660 386 -117632
rect -386 -117928 386 -117900
rect -386 -122162 302 -117928
rect 366 -122162 386 -117928
rect -386 -122190 386 -122162
rect -386 -122458 386 -122430
rect -386 -126692 302 -122458
rect 366 -126692 386 -122458
rect -386 -126720 386 -126692
rect -386 -126988 386 -126960
rect -386 -131222 302 -126988
rect 366 -131222 386 -126988
rect -386 -131250 386 -131222
rect -386 -131518 386 -131490
rect -386 -135752 302 -131518
rect 366 -135752 386 -131518
rect -386 -135780 386 -135752
rect -386 -136048 386 -136020
rect -386 -140282 302 -136048
rect 366 -140282 386 -136048
rect -386 -140310 386 -140282
rect -386 -140578 386 -140550
rect -386 -144812 302 -140578
rect 366 -144812 386 -140578
rect -386 -144840 386 -144812
rect -386 -145108 386 -145080
rect -386 -149342 302 -145108
rect 366 -149342 386 -145108
rect -386 -149370 386 -149342
rect -386 -149638 386 -149610
rect -386 -153872 302 -149638
rect 366 -153872 386 -149638
rect -386 -153900 386 -153872
rect -386 -154168 386 -154140
rect -386 -158402 302 -154168
rect 366 -158402 386 -154168
rect -386 -158430 386 -158402
rect -386 -158698 386 -158670
rect -386 -162932 302 -158698
rect 366 -162932 386 -158698
rect -386 -162960 386 -162932
rect -386 -163228 386 -163200
rect -386 -167462 302 -163228
rect 366 -167462 386 -163228
rect -386 -167490 386 -167462
rect -386 -167758 386 -167730
rect -386 -171992 302 -167758
rect 366 -171992 386 -167758
rect -386 -172020 386 -171992
rect -386 -172288 386 -172260
rect -386 -176522 302 -172288
rect 366 -176522 386 -172288
rect -386 -176550 386 -176522
rect -386 -176818 386 -176790
rect -386 -181052 302 -176818
rect 366 -181052 386 -176818
rect -386 -181080 386 -181052
rect -386 -181348 386 -181320
rect -386 -185582 302 -181348
rect 366 -185582 386 -181348
rect -386 -185610 386 -185582
rect -386 -185878 386 -185850
rect -386 -190112 302 -185878
rect 366 -190112 386 -185878
rect -386 -190140 386 -190112
rect -386 -190408 386 -190380
rect -386 -194642 302 -190408
rect 366 -194642 386 -190408
rect -386 -194670 386 -194642
rect -386 -194938 386 -194910
rect -386 -199172 302 -194938
rect 366 -199172 386 -194938
rect -386 -199200 386 -199172
rect -386 -199468 386 -199440
rect -386 -203702 302 -199468
rect 366 -203702 386 -199468
rect -386 -203730 386 -203702
rect -386 -203998 386 -203970
rect -386 -208232 302 -203998
rect 366 -208232 386 -203998
rect -386 -208260 386 -208232
rect -386 -208528 386 -208500
rect -386 -212762 302 -208528
rect 366 -212762 386 -208528
rect -386 -212790 386 -212762
rect -386 -213058 386 -213030
rect -386 -217292 302 -213058
rect 366 -217292 386 -213058
rect -386 -217320 386 -217292
rect -386 -217588 386 -217560
rect -386 -221822 302 -217588
rect 366 -221822 386 -217588
rect -386 -221850 386 -221822
rect -386 -222118 386 -222090
rect -386 -226352 302 -222118
rect 366 -226352 386 -222118
rect -386 -226380 386 -226352
rect -386 -226648 386 -226620
rect -386 -230882 302 -226648
rect 366 -230882 386 -226648
rect -386 -230910 386 -230882
rect -386 -231178 386 -231150
rect -386 -235412 302 -231178
rect 366 -235412 386 -231178
rect -386 -235440 386 -235412
rect -386 -235708 386 -235680
rect -386 -239942 302 -235708
rect 366 -239942 386 -235708
rect -386 -239970 386 -239942
rect -386 -240238 386 -240210
rect -386 -244472 302 -240238
rect 366 -244472 386 -240238
rect -386 -244500 386 -244472
rect -386 -244768 386 -244740
rect -386 -249002 302 -244768
rect 366 -249002 386 -244768
rect -386 -249030 386 -249002
rect -386 -249298 386 -249270
rect -386 -253532 302 -249298
rect 366 -253532 386 -249298
rect -386 -253560 386 -253532
rect -386 -253828 386 -253800
rect -386 -258062 302 -253828
rect 366 -258062 386 -253828
rect -386 -258090 386 -258062
rect -386 -258358 386 -258330
rect -386 -262592 302 -258358
rect 366 -262592 386 -258358
rect -386 -262620 386 -262592
rect -386 -262888 386 -262860
rect -386 -267122 302 -262888
rect 366 -267122 386 -262888
rect -386 -267150 386 -267122
rect -386 -267418 386 -267390
rect -386 -271652 302 -267418
rect 366 -271652 386 -267418
rect -386 -271680 386 -271652
rect -386 -271948 386 -271920
rect -386 -276182 302 -271948
rect 366 -276182 386 -271948
rect -386 -276210 386 -276182
rect -386 -276478 386 -276450
rect -386 -280712 302 -276478
rect 366 -280712 386 -276478
rect -386 -280740 386 -280712
rect -386 -281008 386 -280980
rect -386 -285242 302 -281008
rect 366 -285242 386 -281008
rect -386 -285270 386 -285242
rect -386 -285538 386 -285510
rect -386 -289772 302 -285538
rect 366 -289772 386 -285538
rect -386 -289800 386 -289772
<< via3 >>
rect 302 285538 366 289772
rect 302 281008 366 285242
rect 302 276478 366 280712
rect 302 271948 366 276182
rect 302 267418 366 271652
rect 302 262888 366 267122
rect 302 258358 366 262592
rect 302 253828 366 258062
rect 302 249298 366 253532
rect 302 244768 366 249002
rect 302 240238 366 244472
rect 302 235708 366 239942
rect 302 231178 366 235412
rect 302 226648 366 230882
rect 302 222118 366 226352
rect 302 217588 366 221822
rect 302 213058 366 217292
rect 302 208528 366 212762
rect 302 203998 366 208232
rect 302 199468 366 203702
rect 302 194938 366 199172
rect 302 190408 366 194642
rect 302 185878 366 190112
rect 302 181348 366 185582
rect 302 176818 366 181052
rect 302 172288 366 176522
rect 302 167758 366 171992
rect 302 163228 366 167462
rect 302 158698 366 162932
rect 302 154168 366 158402
rect 302 149638 366 153872
rect 302 145108 366 149342
rect 302 140578 366 144812
rect 302 136048 366 140282
rect 302 131518 366 135752
rect 302 126988 366 131222
rect 302 122458 366 126692
rect 302 117928 366 122162
rect 302 113398 366 117632
rect 302 108868 366 113102
rect 302 104338 366 108572
rect 302 99808 366 104042
rect 302 95278 366 99512
rect 302 90748 366 94982
rect 302 86218 366 90452
rect 302 81688 366 85922
rect 302 77158 366 81392
rect 302 72628 366 76862
rect 302 68098 366 72332
rect 302 63568 366 67802
rect 302 59038 366 63272
rect 302 54508 366 58742
rect 302 49978 366 54212
rect 302 45448 366 49682
rect 302 40918 366 45152
rect 302 36388 366 40622
rect 302 31858 366 36092
rect 302 27328 366 31562
rect 302 22798 366 27032
rect 302 18268 366 22502
rect 302 13738 366 17972
rect 302 9208 366 13442
rect 302 4678 366 8912
rect 302 148 366 4382
rect 302 -4382 366 -148
rect 302 -8912 366 -4678
rect 302 -13442 366 -9208
rect 302 -17972 366 -13738
rect 302 -22502 366 -18268
rect 302 -27032 366 -22798
rect 302 -31562 366 -27328
rect 302 -36092 366 -31858
rect 302 -40622 366 -36388
rect 302 -45152 366 -40918
rect 302 -49682 366 -45448
rect 302 -54212 366 -49978
rect 302 -58742 366 -54508
rect 302 -63272 366 -59038
rect 302 -67802 366 -63568
rect 302 -72332 366 -68098
rect 302 -76862 366 -72628
rect 302 -81392 366 -77158
rect 302 -85922 366 -81688
rect 302 -90452 366 -86218
rect 302 -94982 366 -90748
rect 302 -99512 366 -95278
rect 302 -104042 366 -99808
rect 302 -108572 366 -104338
rect 302 -113102 366 -108868
rect 302 -117632 366 -113398
rect 302 -122162 366 -117928
rect 302 -126692 366 -122458
rect 302 -131222 366 -126988
rect 302 -135752 366 -131518
rect 302 -140282 366 -136048
rect 302 -144812 366 -140578
rect 302 -149342 366 -145108
rect 302 -153872 366 -149638
rect 302 -158402 366 -154168
rect 302 -162932 366 -158698
rect 302 -167462 366 -163228
rect 302 -171992 366 -167758
rect 302 -176522 366 -172288
rect 302 -181052 366 -176818
rect 302 -185582 366 -181348
rect 302 -190112 366 -185878
rect 302 -194642 366 -190408
rect 302 -199172 366 -194938
rect 302 -203702 366 -199468
rect 302 -208232 366 -203998
rect 302 -212762 366 -208528
rect 302 -217292 366 -213058
rect 302 -221822 366 -217588
rect 302 -226352 366 -222118
rect 302 -230882 366 -226648
rect 302 -235412 366 -231178
rect 302 -239942 366 -235708
rect 302 -244472 366 -240238
rect 302 -249002 366 -244768
rect 302 -253532 366 -249298
rect 302 -258062 366 -253828
rect 302 -262592 366 -258358
rect 302 -267122 366 -262888
rect 302 -271652 366 -267418
rect 302 -276182 366 -271948
rect 302 -280712 366 -276478
rect 302 -285242 366 -281008
rect 302 -289772 366 -285538
<< mimcap >>
rect -346 289720 54 289760
rect -346 285590 -306 289720
rect 14 285590 54 289720
rect -346 285550 54 285590
rect -346 285190 54 285230
rect -346 281060 -306 285190
rect 14 281060 54 285190
rect -346 281020 54 281060
rect -346 280660 54 280700
rect -346 276530 -306 280660
rect 14 276530 54 280660
rect -346 276490 54 276530
rect -346 276130 54 276170
rect -346 272000 -306 276130
rect 14 272000 54 276130
rect -346 271960 54 272000
rect -346 271600 54 271640
rect -346 267470 -306 271600
rect 14 267470 54 271600
rect -346 267430 54 267470
rect -346 267070 54 267110
rect -346 262940 -306 267070
rect 14 262940 54 267070
rect -346 262900 54 262940
rect -346 262540 54 262580
rect -346 258410 -306 262540
rect 14 258410 54 262540
rect -346 258370 54 258410
rect -346 258010 54 258050
rect -346 253880 -306 258010
rect 14 253880 54 258010
rect -346 253840 54 253880
rect -346 253480 54 253520
rect -346 249350 -306 253480
rect 14 249350 54 253480
rect -346 249310 54 249350
rect -346 248950 54 248990
rect -346 244820 -306 248950
rect 14 244820 54 248950
rect -346 244780 54 244820
rect -346 244420 54 244460
rect -346 240290 -306 244420
rect 14 240290 54 244420
rect -346 240250 54 240290
rect -346 239890 54 239930
rect -346 235760 -306 239890
rect 14 235760 54 239890
rect -346 235720 54 235760
rect -346 235360 54 235400
rect -346 231230 -306 235360
rect 14 231230 54 235360
rect -346 231190 54 231230
rect -346 230830 54 230870
rect -346 226700 -306 230830
rect 14 226700 54 230830
rect -346 226660 54 226700
rect -346 226300 54 226340
rect -346 222170 -306 226300
rect 14 222170 54 226300
rect -346 222130 54 222170
rect -346 221770 54 221810
rect -346 217640 -306 221770
rect 14 217640 54 221770
rect -346 217600 54 217640
rect -346 217240 54 217280
rect -346 213110 -306 217240
rect 14 213110 54 217240
rect -346 213070 54 213110
rect -346 212710 54 212750
rect -346 208580 -306 212710
rect 14 208580 54 212710
rect -346 208540 54 208580
rect -346 208180 54 208220
rect -346 204050 -306 208180
rect 14 204050 54 208180
rect -346 204010 54 204050
rect -346 203650 54 203690
rect -346 199520 -306 203650
rect 14 199520 54 203650
rect -346 199480 54 199520
rect -346 199120 54 199160
rect -346 194990 -306 199120
rect 14 194990 54 199120
rect -346 194950 54 194990
rect -346 194590 54 194630
rect -346 190460 -306 194590
rect 14 190460 54 194590
rect -346 190420 54 190460
rect -346 190060 54 190100
rect -346 185930 -306 190060
rect 14 185930 54 190060
rect -346 185890 54 185930
rect -346 185530 54 185570
rect -346 181400 -306 185530
rect 14 181400 54 185530
rect -346 181360 54 181400
rect -346 181000 54 181040
rect -346 176870 -306 181000
rect 14 176870 54 181000
rect -346 176830 54 176870
rect -346 176470 54 176510
rect -346 172340 -306 176470
rect 14 172340 54 176470
rect -346 172300 54 172340
rect -346 171940 54 171980
rect -346 167810 -306 171940
rect 14 167810 54 171940
rect -346 167770 54 167810
rect -346 167410 54 167450
rect -346 163280 -306 167410
rect 14 163280 54 167410
rect -346 163240 54 163280
rect -346 162880 54 162920
rect -346 158750 -306 162880
rect 14 158750 54 162880
rect -346 158710 54 158750
rect -346 158350 54 158390
rect -346 154220 -306 158350
rect 14 154220 54 158350
rect -346 154180 54 154220
rect -346 153820 54 153860
rect -346 149690 -306 153820
rect 14 149690 54 153820
rect -346 149650 54 149690
rect -346 149290 54 149330
rect -346 145160 -306 149290
rect 14 145160 54 149290
rect -346 145120 54 145160
rect -346 144760 54 144800
rect -346 140630 -306 144760
rect 14 140630 54 144760
rect -346 140590 54 140630
rect -346 140230 54 140270
rect -346 136100 -306 140230
rect 14 136100 54 140230
rect -346 136060 54 136100
rect -346 135700 54 135740
rect -346 131570 -306 135700
rect 14 131570 54 135700
rect -346 131530 54 131570
rect -346 131170 54 131210
rect -346 127040 -306 131170
rect 14 127040 54 131170
rect -346 127000 54 127040
rect -346 126640 54 126680
rect -346 122510 -306 126640
rect 14 122510 54 126640
rect -346 122470 54 122510
rect -346 122110 54 122150
rect -346 117980 -306 122110
rect 14 117980 54 122110
rect -346 117940 54 117980
rect -346 117580 54 117620
rect -346 113450 -306 117580
rect 14 113450 54 117580
rect -346 113410 54 113450
rect -346 113050 54 113090
rect -346 108920 -306 113050
rect 14 108920 54 113050
rect -346 108880 54 108920
rect -346 108520 54 108560
rect -346 104390 -306 108520
rect 14 104390 54 108520
rect -346 104350 54 104390
rect -346 103990 54 104030
rect -346 99860 -306 103990
rect 14 99860 54 103990
rect -346 99820 54 99860
rect -346 99460 54 99500
rect -346 95330 -306 99460
rect 14 95330 54 99460
rect -346 95290 54 95330
rect -346 94930 54 94970
rect -346 90800 -306 94930
rect 14 90800 54 94930
rect -346 90760 54 90800
rect -346 90400 54 90440
rect -346 86270 -306 90400
rect 14 86270 54 90400
rect -346 86230 54 86270
rect -346 85870 54 85910
rect -346 81740 -306 85870
rect 14 81740 54 85870
rect -346 81700 54 81740
rect -346 81340 54 81380
rect -346 77210 -306 81340
rect 14 77210 54 81340
rect -346 77170 54 77210
rect -346 76810 54 76850
rect -346 72680 -306 76810
rect 14 72680 54 76810
rect -346 72640 54 72680
rect -346 72280 54 72320
rect -346 68150 -306 72280
rect 14 68150 54 72280
rect -346 68110 54 68150
rect -346 67750 54 67790
rect -346 63620 -306 67750
rect 14 63620 54 67750
rect -346 63580 54 63620
rect -346 63220 54 63260
rect -346 59090 -306 63220
rect 14 59090 54 63220
rect -346 59050 54 59090
rect -346 58690 54 58730
rect -346 54560 -306 58690
rect 14 54560 54 58690
rect -346 54520 54 54560
rect -346 54160 54 54200
rect -346 50030 -306 54160
rect 14 50030 54 54160
rect -346 49990 54 50030
rect -346 49630 54 49670
rect -346 45500 -306 49630
rect 14 45500 54 49630
rect -346 45460 54 45500
rect -346 45100 54 45140
rect -346 40970 -306 45100
rect 14 40970 54 45100
rect -346 40930 54 40970
rect -346 40570 54 40610
rect -346 36440 -306 40570
rect 14 36440 54 40570
rect -346 36400 54 36440
rect -346 36040 54 36080
rect -346 31910 -306 36040
rect 14 31910 54 36040
rect -346 31870 54 31910
rect -346 31510 54 31550
rect -346 27380 -306 31510
rect 14 27380 54 31510
rect -346 27340 54 27380
rect -346 26980 54 27020
rect -346 22850 -306 26980
rect 14 22850 54 26980
rect -346 22810 54 22850
rect -346 22450 54 22490
rect -346 18320 -306 22450
rect 14 18320 54 22450
rect -346 18280 54 18320
rect -346 17920 54 17960
rect -346 13790 -306 17920
rect 14 13790 54 17920
rect -346 13750 54 13790
rect -346 13390 54 13430
rect -346 9260 -306 13390
rect 14 9260 54 13390
rect -346 9220 54 9260
rect -346 8860 54 8900
rect -346 4730 -306 8860
rect 14 4730 54 8860
rect -346 4690 54 4730
rect -346 4330 54 4370
rect -346 200 -306 4330
rect 14 200 54 4330
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -4330 -306 -200
rect 14 -4330 54 -200
rect -346 -4370 54 -4330
rect -346 -4730 54 -4690
rect -346 -8860 -306 -4730
rect 14 -8860 54 -4730
rect -346 -8900 54 -8860
rect -346 -9260 54 -9220
rect -346 -13390 -306 -9260
rect 14 -13390 54 -9260
rect -346 -13430 54 -13390
rect -346 -13790 54 -13750
rect -346 -17920 -306 -13790
rect 14 -17920 54 -13790
rect -346 -17960 54 -17920
rect -346 -18320 54 -18280
rect -346 -22450 -306 -18320
rect 14 -22450 54 -18320
rect -346 -22490 54 -22450
rect -346 -22850 54 -22810
rect -346 -26980 -306 -22850
rect 14 -26980 54 -22850
rect -346 -27020 54 -26980
rect -346 -27380 54 -27340
rect -346 -31510 -306 -27380
rect 14 -31510 54 -27380
rect -346 -31550 54 -31510
rect -346 -31910 54 -31870
rect -346 -36040 -306 -31910
rect 14 -36040 54 -31910
rect -346 -36080 54 -36040
rect -346 -36440 54 -36400
rect -346 -40570 -306 -36440
rect 14 -40570 54 -36440
rect -346 -40610 54 -40570
rect -346 -40970 54 -40930
rect -346 -45100 -306 -40970
rect 14 -45100 54 -40970
rect -346 -45140 54 -45100
rect -346 -45500 54 -45460
rect -346 -49630 -306 -45500
rect 14 -49630 54 -45500
rect -346 -49670 54 -49630
rect -346 -50030 54 -49990
rect -346 -54160 -306 -50030
rect 14 -54160 54 -50030
rect -346 -54200 54 -54160
rect -346 -54560 54 -54520
rect -346 -58690 -306 -54560
rect 14 -58690 54 -54560
rect -346 -58730 54 -58690
rect -346 -59090 54 -59050
rect -346 -63220 -306 -59090
rect 14 -63220 54 -59090
rect -346 -63260 54 -63220
rect -346 -63620 54 -63580
rect -346 -67750 -306 -63620
rect 14 -67750 54 -63620
rect -346 -67790 54 -67750
rect -346 -68150 54 -68110
rect -346 -72280 -306 -68150
rect 14 -72280 54 -68150
rect -346 -72320 54 -72280
rect -346 -72680 54 -72640
rect -346 -76810 -306 -72680
rect 14 -76810 54 -72680
rect -346 -76850 54 -76810
rect -346 -77210 54 -77170
rect -346 -81340 -306 -77210
rect 14 -81340 54 -77210
rect -346 -81380 54 -81340
rect -346 -81740 54 -81700
rect -346 -85870 -306 -81740
rect 14 -85870 54 -81740
rect -346 -85910 54 -85870
rect -346 -86270 54 -86230
rect -346 -90400 -306 -86270
rect 14 -90400 54 -86270
rect -346 -90440 54 -90400
rect -346 -90800 54 -90760
rect -346 -94930 -306 -90800
rect 14 -94930 54 -90800
rect -346 -94970 54 -94930
rect -346 -95330 54 -95290
rect -346 -99460 -306 -95330
rect 14 -99460 54 -95330
rect -346 -99500 54 -99460
rect -346 -99860 54 -99820
rect -346 -103990 -306 -99860
rect 14 -103990 54 -99860
rect -346 -104030 54 -103990
rect -346 -104390 54 -104350
rect -346 -108520 -306 -104390
rect 14 -108520 54 -104390
rect -346 -108560 54 -108520
rect -346 -108920 54 -108880
rect -346 -113050 -306 -108920
rect 14 -113050 54 -108920
rect -346 -113090 54 -113050
rect -346 -113450 54 -113410
rect -346 -117580 -306 -113450
rect 14 -117580 54 -113450
rect -346 -117620 54 -117580
rect -346 -117980 54 -117940
rect -346 -122110 -306 -117980
rect 14 -122110 54 -117980
rect -346 -122150 54 -122110
rect -346 -122510 54 -122470
rect -346 -126640 -306 -122510
rect 14 -126640 54 -122510
rect -346 -126680 54 -126640
rect -346 -127040 54 -127000
rect -346 -131170 -306 -127040
rect 14 -131170 54 -127040
rect -346 -131210 54 -131170
rect -346 -131570 54 -131530
rect -346 -135700 -306 -131570
rect 14 -135700 54 -131570
rect -346 -135740 54 -135700
rect -346 -136100 54 -136060
rect -346 -140230 -306 -136100
rect 14 -140230 54 -136100
rect -346 -140270 54 -140230
rect -346 -140630 54 -140590
rect -346 -144760 -306 -140630
rect 14 -144760 54 -140630
rect -346 -144800 54 -144760
rect -346 -145160 54 -145120
rect -346 -149290 -306 -145160
rect 14 -149290 54 -145160
rect -346 -149330 54 -149290
rect -346 -149690 54 -149650
rect -346 -153820 -306 -149690
rect 14 -153820 54 -149690
rect -346 -153860 54 -153820
rect -346 -154220 54 -154180
rect -346 -158350 -306 -154220
rect 14 -158350 54 -154220
rect -346 -158390 54 -158350
rect -346 -158750 54 -158710
rect -346 -162880 -306 -158750
rect 14 -162880 54 -158750
rect -346 -162920 54 -162880
rect -346 -163280 54 -163240
rect -346 -167410 -306 -163280
rect 14 -167410 54 -163280
rect -346 -167450 54 -167410
rect -346 -167810 54 -167770
rect -346 -171940 -306 -167810
rect 14 -171940 54 -167810
rect -346 -171980 54 -171940
rect -346 -172340 54 -172300
rect -346 -176470 -306 -172340
rect 14 -176470 54 -172340
rect -346 -176510 54 -176470
rect -346 -176870 54 -176830
rect -346 -181000 -306 -176870
rect 14 -181000 54 -176870
rect -346 -181040 54 -181000
rect -346 -181400 54 -181360
rect -346 -185530 -306 -181400
rect 14 -185530 54 -181400
rect -346 -185570 54 -185530
rect -346 -185930 54 -185890
rect -346 -190060 -306 -185930
rect 14 -190060 54 -185930
rect -346 -190100 54 -190060
rect -346 -190460 54 -190420
rect -346 -194590 -306 -190460
rect 14 -194590 54 -190460
rect -346 -194630 54 -194590
rect -346 -194990 54 -194950
rect -346 -199120 -306 -194990
rect 14 -199120 54 -194990
rect -346 -199160 54 -199120
rect -346 -199520 54 -199480
rect -346 -203650 -306 -199520
rect 14 -203650 54 -199520
rect -346 -203690 54 -203650
rect -346 -204050 54 -204010
rect -346 -208180 -306 -204050
rect 14 -208180 54 -204050
rect -346 -208220 54 -208180
rect -346 -208580 54 -208540
rect -346 -212710 -306 -208580
rect 14 -212710 54 -208580
rect -346 -212750 54 -212710
rect -346 -213110 54 -213070
rect -346 -217240 -306 -213110
rect 14 -217240 54 -213110
rect -346 -217280 54 -217240
rect -346 -217640 54 -217600
rect -346 -221770 -306 -217640
rect 14 -221770 54 -217640
rect -346 -221810 54 -221770
rect -346 -222170 54 -222130
rect -346 -226300 -306 -222170
rect 14 -226300 54 -222170
rect -346 -226340 54 -226300
rect -346 -226700 54 -226660
rect -346 -230830 -306 -226700
rect 14 -230830 54 -226700
rect -346 -230870 54 -230830
rect -346 -231230 54 -231190
rect -346 -235360 -306 -231230
rect 14 -235360 54 -231230
rect -346 -235400 54 -235360
rect -346 -235760 54 -235720
rect -346 -239890 -306 -235760
rect 14 -239890 54 -235760
rect -346 -239930 54 -239890
rect -346 -240290 54 -240250
rect -346 -244420 -306 -240290
rect 14 -244420 54 -240290
rect -346 -244460 54 -244420
rect -346 -244820 54 -244780
rect -346 -248950 -306 -244820
rect 14 -248950 54 -244820
rect -346 -248990 54 -248950
rect -346 -249350 54 -249310
rect -346 -253480 -306 -249350
rect 14 -253480 54 -249350
rect -346 -253520 54 -253480
rect -346 -253880 54 -253840
rect -346 -258010 -306 -253880
rect 14 -258010 54 -253880
rect -346 -258050 54 -258010
rect -346 -258410 54 -258370
rect -346 -262540 -306 -258410
rect 14 -262540 54 -258410
rect -346 -262580 54 -262540
rect -346 -262940 54 -262900
rect -346 -267070 -306 -262940
rect 14 -267070 54 -262940
rect -346 -267110 54 -267070
rect -346 -267470 54 -267430
rect -346 -271600 -306 -267470
rect 14 -271600 54 -267470
rect -346 -271640 54 -271600
rect -346 -272000 54 -271960
rect -346 -276130 -306 -272000
rect 14 -276130 54 -272000
rect -346 -276170 54 -276130
rect -346 -276530 54 -276490
rect -346 -280660 -306 -276530
rect 14 -280660 54 -276530
rect -346 -280700 54 -280660
rect -346 -281060 54 -281020
rect -346 -285190 -306 -281060
rect 14 -285190 54 -281060
rect -346 -285230 54 -285190
rect -346 -285590 54 -285550
rect -346 -289720 -306 -285590
rect 14 -289720 54 -285590
rect -346 -289760 54 -289720
<< mimcapcontact >>
rect -306 285590 14 289720
rect -306 281060 14 285190
rect -306 276530 14 280660
rect -306 272000 14 276130
rect -306 267470 14 271600
rect -306 262940 14 267070
rect -306 258410 14 262540
rect -306 253880 14 258010
rect -306 249350 14 253480
rect -306 244820 14 248950
rect -306 240290 14 244420
rect -306 235760 14 239890
rect -306 231230 14 235360
rect -306 226700 14 230830
rect -306 222170 14 226300
rect -306 217640 14 221770
rect -306 213110 14 217240
rect -306 208580 14 212710
rect -306 204050 14 208180
rect -306 199520 14 203650
rect -306 194990 14 199120
rect -306 190460 14 194590
rect -306 185930 14 190060
rect -306 181400 14 185530
rect -306 176870 14 181000
rect -306 172340 14 176470
rect -306 167810 14 171940
rect -306 163280 14 167410
rect -306 158750 14 162880
rect -306 154220 14 158350
rect -306 149690 14 153820
rect -306 145160 14 149290
rect -306 140630 14 144760
rect -306 136100 14 140230
rect -306 131570 14 135700
rect -306 127040 14 131170
rect -306 122510 14 126640
rect -306 117980 14 122110
rect -306 113450 14 117580
rect -306 108920 14 113050
rect -306 104390 14 108520
rect -306 99860 14 103990
rect -306 95330 14 99460
rect -306 90800 14 94930
rect -306 86270 14 90400
rect -306 81740 14 85870
rect -306 77210 14 81340
rect -306 72680 14 76810
rect -306 68150 14 72280
rect -306 63620 14 67750
rect -306 59090 14 63220
rect -306 54560 14 58690
rect -306 50030 14 54160
rect -306 45500 14 49630
rect -306 40970 14 45100
rect -306 36440 14 40570
rect -306 31910 14 36040
rect -306 27380 14 31510
rect -306 22850 14 26980
rect -306 18320 14 22450
rect -306 13790 14 17920
rect -306 9260 14 13390
rect -306 4730 14 8860
rect -306 200 14 4330
rect -306 -4330 14 -200
rect -306 -8860 14 -4730
rect -306 -13390 14 -9260
rect -306 -17920 14 -13790
rect -306 -22450 14 -18320
rect -306 -26980 14 -22850
rect -306 -31510 14 -27380
rect -306 -36040 14 -31910
rect -306 -40570 14 -36440
rect -306 -45100 14 -40970
rect -306 -49630 14 -45500
rect -306 -54160 14 -50030
rect -306 -58690 14 -54560
rect -306 -63220 14 -59090
rect -306 -67750 14 -63620
rect -306 -72280 14 -68150
rect -306 -76810 14 -72680
rect -306 -81340 14 -77210
rect -306 -85870 14 -81740
rect -306 -90400 14 -86270
rect -306 -94930 14 -90800
rect -306 -99460 14 -95330
rect -306 -103990 14 -99860
rect -306 -108520 14 -104390
rect -306 -113050 14 -108920
rect -306 -117580 14 -113450
rect -306 -122110 14 -117980
rect -306 -126640 14 -122510
rect -306 -131170 14 -127040
rect -306 -135700 14 -131570
rect -306 -140230 14 -136100
rect -306 -144760 14 -140630
rect -306 -149290 14 -145160
rect -306 -153820 14 -149690
rect -306 -158350 14 -154220
rect -306 -162880 14 -158750
rect -306 -167410 14 -163280
rect -306 -171940 14 -167810
rect -306 -176470 14 -172340
rect -306 -181000 14 -176870
rect -306 -185530 14 -181400
rect -306 -190060 14 -185930
rect -306 -194590 14 -190460
rect -306 -199120 14 -194990
rect -306 -203650 14 -199520
rect -306 -208180 14 -204050
rect -306 -212710 14 -208580
rect -306 -217240 14 -213110
rect -306 -221770 14 -217640
rect -306 -226300 14 -222170
rect -306 -230830 14 -226700
rect -306 -235360 14 -231230
rect -306 -239890 14 -235760
rect -306 -244420 14 -240290
rect -306 -248950 14 -244820
rect -306 -253480 14 -249350
rect -306 -258010 14 -253880
rect -306 -262540 14 -258410
rect -306 -267070 14 -262940
rect -306 -271600 14 -267470
rect -306 -276130 14 -272000
rect -306 -280660 14 -276530
rect -306 -285190 14 -281060
rect -306 -289720 14 -285590
<< metal4 >>
rect -198 289721 -94 289920
rect 282 289772 386 289920
rect -307 289720 15 289721
rect -307 285590 -306 289720
rect 14 285590 15 289720
rect -307 285589 15 285590
rect -198 285191 -94 285589
rect 282 285538 302 289772
rect 366 285538 386 289772
rect 282 285242 386 285538
rect -307 285190 15 285191
rect -307 281060 -306 285190
rect 14 281060 15 285190
rect -307 281059 15 281060
rect -198 280661 -94 281059
rect 282 281008 302 285242
rect 366 281008 386 285242
rect 282 280712 386 281008
rect -307 280660 15 280661
rect -307 276530 -306 280660
rect 14 276530 15 280660
rect -307 276529 15 276530
rect -198 276131 -94 276529
rect 282 276478 302 280712
rect 366 276478 386 280712
rect 282 276182 386 276478
rect -307 276130 15 276131
rect -307 272000 -306 276130
rect 14 272000 15 276130
rect -307 271999 15 272000
rect -198 271601 -94 271999
rect 282 271948 302 276182
rect 366 271948 386 276182
rect 282 271652 386 271948
rect -307 271600 15 271601
rect -307 267470 -306 271600
rect 14 267470 15 271600
rect -307 267469 15 267470
rect -198 267071 -94 267469
rect 282 267418 302 271652
rect 366 267418 386 271652
rect 282 267122 386 267418
rect -307 267070 15 267071
rect -307 262940 -306 267070
rect 14 262940 15 267070
rect -307 262939 15 262940
rect -198 262541 -94 262939
rect 282 262888 302 267122
rect 366 262888 386 267122
rect 282 262592 386 262888
rect -307 262540 15 262541
rect -307 258410 -306 262540
rect 14 258410 15 262540
rect -307 258409 15 258410
rect -198 258011 -94 258409
rect 282 258358 302 262592
rect 366 258358 386 262592
rect 282 258062 386 258358
rect -307 258010 15 258011
rect -307 253880 -306 258010
rect 14 253880 15 258010
rect -307 253879 15 253880
rect -198 253481 -94 253879
rect 282 253828 302 258062
rect 366 253828 386 258062
rect 282 253532 386 253828
rect -307 253480 15 253481
rect -307 249350 -306 253480
rect 14 249350 15 253480
rect -307 249349 15 249350
rect -198 248951 -94 249349
rect 282 249298 302 253532
rect 366 249298 386 253532
rect 282 249002 386 249298
rect -307 248950 15 248951
rect -307 244820 -306 248950
rect 14 244820 15 248950
rect -307 244819 15 244820
rect -198 244421 -94 244819
rect 282 244768 302 249002
rect 366 244768 386 249002
rect 282 244472 386 244768
rect -307 244420 15 244421
rect -307 240290 -306 244420
rect 14 240290 15 244420
rect -307 240289 15 240290
rect -198 239891 -94 240289
rect 282 240238 302 244472
rect 366 240238 386 244472
rect 282 239942 386 240238
rect -307 239890 15 239891
rect -307 235760 -306 239890
rect 14 235760 15 239890
rect -307 235759 15 235760
rect -198 235361 -94 235759
rect 282 235708 302 239942
rect 366 235708 386 239942
rect 282 235412 386 235708
rect -307 235360 15 235361
rect -307 231230 -306 235360
rect 14 231230 15 235360
rect -307 231229 15 231230
rect -198 230831 -94 231229
rect 282 231178 302 235412
rect 366 231178 386 235412
rect 282 230882 386 231178
rect -307 230830 15 230831
rect -307 226700 -306 230830
rect 14 226700 15 230830
rect -307 226699 15 226700
rect -198 226301 -94 226699
rect 282 226648 302 230882
rect 366 226648 386 230882
rect 282 226352 386 226648
rect -307 226300 15 226301
rect -307 222170 -306 226300
rect 14 222170 15 226300
rect -307 222169 15 222170
rect -198 221771 -94 222169
rect 282 222118 302 226352
rect 366 222118 386 226352
rect 282 221822 386 222118
rect -307 221770 15 221771
rect -307 217640 -306 221770
rect 14 217640 15 221770
rect -307 217639 15 217640
rect -198 217241 -94 217639
rect 282 217588 302 221822
rect 366 217588 386 221822
rect 282 217292 386 217588
rect -307 217240 15 217241
rect -307 213110 -306 217240
rect 14 213110 15 217240
rect -307 213109 15 213110
rect -198 212711 -94 213109
rect 282 213058 302 217292
rect 366 213058 386 217292
rect 282 212762 386 213058
rect -307 212710 15 212711
rect -307 208580 -306 212710
rect 14 208580 15 212710
rect -307 208579 15 208580
rect -198 208181 -94 208579
rect 282 208528 302 212762
rect 366 208528 386 212762
rect 282 208232 386 208528
rect -307 208180 15 208181
rect -307 204050 -306 208180
rect 14 204050 15 208180
rect -307 204049 15 204050
rect -198 203651 -94 204049
rect 282 203998 302 208232
rect 366 203998 386 208232
rect 282 203702 386 203998
rect -307 203650 15 203651
rect -307 199520 -306 203650
rect 14 199520 15 203650
rect -307 199519 15 199520
rect -198 199121 -94 199519
rect 282 199468 302 203702
rect 366 199468 386 203702
rect 282 199172 386 199468
rect -307 199120 15 199121
rect -307 194990 -306 199120
rect 14 194990 15 199120
rect -307 194989 15 194990
rect -198 194591 -94 194989
rect 282 194938 302 199172
rect 366 194938 386 199172
rect 282 194642 386 194938
rect -307 194590 15 194591
rect -307 190460 -306 194590
rect 14 190460 15 194590
rect -307 190459 15 190460
rect -198 190061 -94 190459
rect 282 190408 302 194642
rect 366 190408 386 194642
rect 282 190112 386 190408
rect -307 190060 15 190061
rect -307 185930 -306 190060
rect 14 185930 15 190060
rect -307 185929 15 185930
rect -198 185531 -94 185929
rect 282 185878 302 190112
rect 366 185878 386 190112
rect 282 185582 386 185878
rect -307 185530 15 185531
rect -307 181400 -306 185530
rect 14 181400 15 185530
rect -307 181399 15 181400
rect -198 181001 -94 181399
rect 282 181348 302 185582
rect 366 181348 386 185582
rect 282 181052 386 181348
rect -307 181000 15 181001
rect -307 176870 -306 181000
rect 14 176870 15 181000
rect -307 176869 15 176870
rect -198 176471 -94 176869
rect 282 176818 302 181052
rect 366 176818 386 181052
rect 282 176522 386 176818
rect -307 176470 15 176471
rect -307 172340 -306 176470
rect 14 172340 15 176470
rect -307 172339 15 172340
rect -198 171941 -94 172339
rect 282 172288 302 176522
rect 366 172288 386 176522
rect 282 171992 386 172288
rect -307 171940 15 171941
rect -307 167810 -306 171940
rect 14 167810 15 171940
rect -307 167809 15 167810
rect -198 167411 -94 167809
rect 282 167758 302 171992
rect 366 167758 386 171992
rect 282 167462 386 167758
rect -307 167410 15 167411
rect -307 163280 -306 167410
rect 14 163280 15 167410
rect -307 163279 15 163280
rect -198 162881 -94 163279
rect 282 163228 302 167462
rect 366 163228 386 167462
rect 282 162932 386 163228
rect -307 162880 15 162881
rect -307 158750 -306 162880
rect 14 158750 15 162880
rect -307 158749 15 158750
rect -198 158351 -94 158749
rect 282 158698 302 162932
rect 366 158698 386 162932
rect 282 158402 386 158698
rect -307 158350 15 158351
rect -307 154220 -306 158350
rect 14 154220 15 158350
rect -307 154219 15 154220
rect -198 153821 -94 154219
rect 282 154168 302 158402
rect 366 154168 386 158402
rect 282 153872 386 154168
rect -307 153820 15 153821
rect -307 149690 -306 153820
rect 14 149690 15 153820
rect -307 149689 15 149690
rect -198 149291 -94 149689
rect 282 149638 302 153872
rect 366 149638 386 153872
rect 282 149342 386 149638
rect -307 149290 15 149291
rect -307 145160 -306 149290
rect 14 145160 15 149290
rect -307 145159 15 145160
rect -198 144761 -94 145159
rect 282 145108 302 149342
rect 366 145108 386 149342
rect 282 144812 386 145108
rect -307 144760 15 144761
rect -307 140630 -306 144760
rect 14 140630 15 144760
rect -307 140629 15 140630
rect -198 140231 -94 140629
rect 282 140578 302 144812
rect 366 140578 386 144812
rect 282 140282 386 140578
rect -307 140230 15 140231
rect -307 136100 -306 140230
rect 14 136100 15 140230
rect -307 136099 15 136100
rect -198 135701 -94 136099
rect 282 136048 302 140282
rect 366 136048 386 140282
rect 282 135752 386 136048
rect -307 135700 15 135701
rect -307 131570 -306 135700
rect 14 131570 15 135700
rect -307 131569 15 131570
rect -198 131171 -94 131569
rect 282 131518 302 135752
rect 366 131518 386 135752
rect 282 131222 386 131518
rect -307 131170 15 131171
rect -307 127040 -306 131170
rect 14 127040 15 131170
rect -307 127039 15 127040
rect -198 126641 -94 127039
rect 282 126988 302 131222
rect 366 126988 386 131222
rect 282 126692 386 126988
rect -307 126640 15 126641
rect -307 122510 -306 126640
rect 14 122510 15 126640
rect -307 122509 15 122510
rect -198 122111 -94 122509
rect 282 122458 302 126692
rect 366 122458 386 126692
rect 282 122162 386 122458
rect -307 122110 15 122111
rect -307 117980 -306 122110
rect 14 117980 15 122110
rect -307 117979 15 117980
rect -198 117581 -94 117979
rect 282 117928 302 122162
rect 366 117928 386 122162
rect 282 117632 386 117928
rect -307 117580 15 117581
rect -307 113450 -306 117580
rect 14 113450 15 117580
rect -307 113449 15 113450
rect -198 113051 -94 113449
rect 282 113398 302 117632
rect 366 113398 386 117632
rect 282 113102 386 113398
rect -307 113050 15 113051
rect -307 108920 -306 113050
rect 14 108920 15 113050
rect -307 108919 15 108920
rect -198 108521 -94 108919
rect 282 108868 302 113102
rect 366 108868 386 113102
rect 282 108572 386 108868
rect -307 108520 15 108521
rect -307 104390 -306 108520
rect 14 104390 15 108520
rect -307 104389 15 104390
rect -198 103991 -94 104389
rect 282 104338 302 108572
rect 366 104338 386 108572
rect 282 104042 386 104338
rect -307 103990 15 103991
rect -307 99860 -306 103990
rect 14 99860 15 103990
rect -307 99859 15 99860
rect -198 99461 -94 99859
rect 282 99808 302 104042
rect 366 99808 386 104042
rect 282 99512 386 99808
rect -307 99460 15 99461
rect -307 95330 -306 99460
rect 14 95330 15 99460
rect -307 95329 15 95330
rect -198 94931 -94 95329
rect 282 95278 302 99512
rect 366 95278 386 99512
rect 282 94982 386 95278
rect -307 94930 15 94931
rect -307 90800 -306 94930
rect 14 90800 15 94930
rect -307 90799 15 90800
rect -198 90401 -94 90799
rect 282 90748 302 94982
rect 366 90748 386 94982
rect 282 90452 386 90748
rect -307 90400 15 90401
rect -307 86270 -306 90400
rect 14 86270 15 90400
rect -307 86269 15 86270
rect -198 85871 -94 86269
rect 282 86218 302 90452
rect 366 86218 386 90452
rect 282 85922 386 86218
rect -307 85870 15 85871
rect -307 81740 -306 85870
rect 14 81740 15 85870
rect -307 81739 15 81740
rect -198 81341 -94 81739
rect 282 81688 302 85922
rect 366 81688 386 85922
rect 282 81392 386 81688
rect -307 81340 15 81341
rect -307 77210 -306 81340
rect 14 77210 15 81340
rect -307 77209 15 77210
rect -198 76811 -94 77209
rect 282 77158 302 81392
rect 366 77158 386 81392
rect 282 76862 386 77158
rect -307 76810 15 76811
rect -307 72680 -306 76810
rect 14 72680 15 76810
rect -307 72679 15 72680
rect -198 72281 -94 72679
rect 282 72628 302 76862
rect 366 72628 386 76862
rect 282 72332 386 72628
rect -307 72280 15 72281
rect -307 68150 -306 72280
rect 14 68150 15 72280
rect -307 68149 15 68150
rect -198 67751 -94 68149
rect 282 68098 302 72332
rect 366 68098 386 72332
rect 282 67802 386 68098
rect -307 67750 15 67751
rect -307 63620 -306 67750
rect 14 63620 15 67750
rect -307 63619 15 63620
rect -198 63221 -94 63619
rect 282 63568 302 67802
rect 366 63568 386 67802
rect 282 63272 386 63568
rect -307 63220 15 63221
rect -307 59090 -306 63220
rect 14 59090 15 63220
rect -307 59089 15 59090
rect -198 58691 -94 59089
rect 282 59038 302 63272
rect 366 59038 386 63272
rect 282 58742 386 59038
rect -307 58690 15 58691
rect -307 54560 -306 58690
rect 14 54560 15 58690
rect -307 54559 15 54560
rect -198 54161 -94 54559
rect 282 54508 302 58742
rect 366 54508 386 58742
rect 282 54212 386 54508
rect -307 54160 15 54161
rect -307 50030 -306 54160
rect 14 50030 15 54160
rect -307 50029 15 50030
rect -198 49631 -94 50029
rect 282 49978 302 54212
rect 366 49978 386 54212
rect 282 49682 386 49978
rect -307 49630 15 49631
rect -307 45500 -306 49630
rect 14 45500 15 49630
rect -307 45499 15 45500
rect -198 45101 -94 45499
rect 282 45448 302 49682
rect 366 45448 386 49682
rect 282 45152 386 45448
rect -307 45100 15 45101
rect -307 40970 -306 45100
rect 14 40970 15 45100
rect -307 40969 15 40970
rect -198 40571 -94 40969
rect 282 40918 302 45152
rect 366 40918 386 45152
rect 282 40622 386 40918
rect -307 40570 15 40571
rect -307 36440 -306 40570
rect 14 36440 15 40570
rect -307 36439 15 36440
rect -198 36041 -94 36439
rect 282 36388 302 40622
rect 366 36388 386 40622
rect 282 36092 386 36388
rect -307 36040 15 36041
rect -307 31910 -306 36040
rect 14 31910 15 36040
rect -307 31909 15 31910
rect -198 31511 -94 31909
rect 282 31858 302 36092
rect 366 31858 386 36092
rect 282 31562 386 31858
rect -307 31510 15 31511
rect -307 27380 -306 31510
rect 14 27380 15 31510
rect -307 27379 15 27380
rect -198 26981 -94 27379
rect 282 27328 302 31562
rect 366 27328 386 31562
rect 282 27032 386 27328
rect -307 26980 15 26981
rect -307 22850 -306 26980
rect 14 22850 15 26980
rect -307 22849 15 22850
rect -198 22451 -94 22849
rect 282 22798 302 27032
rect 366 22798 386 27032
rect 282 22502 386 22798
rect -307 22450 15 22451
rect -307 18320 -306 22450
rect 14 18320 15 22450
rect -307 18319 15 18320
rect -198 17921 -94 18319
rect 282 18268 302 22502
rect 366 18268 386 22502
rect 282 17972 386 18268
rect -307 17920 15 17921
rect -307 13790 -306 17920
rect 14 13790 15 17920
rect -307 13789 15 13790
rect -198 13391 -94 13789
rect 282 13738 302 17972
rect 366 13738 386 17972
rect 282 13442 386 13738
rect -307 13390 15 13391
rect -307 9260 -306 13390
rect 14 9260 15 13390
rect -307 9259 15 9260
rect -198 8861 -94 9259
rect 282 9208 302 13442
rect 366 9208 386 13442
rect 282 8912 386 9208
rect -307 8860 15 8861
rect -307 4730 -306 8860
rect 14 4730 15 8860
rect -307 4729 15 4730
rect -198 4331 -94 4729
rect 282 4678 302 8912
rect 366 4678 386 8912
rect 282 4382 386 4678
rect -307 4330 15 4331
rect -307 200 -306 4330
rect 14 200 15 4330
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 4382
rect 366 148 386 4382
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -4330 -306 -200
rect 14 -4330 15 -200
rect -307 -4331 15 -4330
rect -198 -4729 -94 -4331
rect 282 -4382 302 -148
rect 366 -4382 386 -148
rect 282 -4678 386 -4382
rect -307 -4730 15 -4729
rect -307 -8860 -306 -4730
rect 14 -8860 15 -4730
rect -307 -8861 15 -8860
rect -198 -9259 -94 -8861
rect 282 -8912 302 -4678
rect 366 -8912 386 -4678
rect 282 -9208 386 -8912
rect -307 -9260 15 -9259
rect -307 -13390 -306 -9260
rect 14 -13390 15 -9260
rect -307 -13391 15 -13390
rect -198 -13789 -94 -13391
rect 282 -13442 302 -9208
rect 366 -13442 386 -9208
rect 282 -13738 386 -13442
rect -307 -13790 15 -13789
rect -307 -17920 -306 -13790
rect 14 -17920 15 -13790
rect -307 -17921 15 -17920
rect -198 -18319 -94 -17921
rect 282 -17972 302 -13738
rect 366 -17972 386 -13738
rect 282 -18268 386 -17972
rect -307 -18320 15 -18319
rect -307 -22450 -306 -18320
rect 14 -22450 15 -18320
rect -307 -22451 15 -22450
rect -198 -22849 -94 -22451
rect 282 -22502 302 -18268
rect 366 -22502 386 -18268
rect 282 -22798 386 -22502
rect -307 -22850 15 -22849
rect -307 -26980 -306 -22850
rect 14 -26980 15 -22850
rect -307 -26981 15 -26980
rect -198 -27379 -94 -26981
rect 282 -27032 302 -22798
rect 366 -27032 386 -22798
rect 282 -27328 386 -27032
rect -307 -27380 15 -27379
rect -307 -31510 -306 -27380
rect 14 -31510 15 -27380
rect -307 -31511 15 -31510
rect -198 -31909 -94 -31511
rect 282 -31562 302 -27328
rect 366 -31562 386 -27328
rect 282 -31858 386 -31562
rect -307 -31910 15 -31909
rect -307 -36040 -306 -31910
rect 14 -36040 15 -31910
rect -307 -36041 15 -36040
rect -198 -36439 -94 -36041
rect 282 -36092 302 -31858
rect 366 -36092 386 -31858
rect 282 -36388 386 -36092
rect -307 -36440 15 -36439
rect -307 -40570 -306 -36440
rect 14 -40570 15 -36440
rect -307 -40571 15 -40570
rect -198 -40969 -94 -40571
rect 282 -40622 302 -36388
rect 366 -40622 386 -36388
rect 282 -40918 386 -40622
rect -307 -40970 15 -40969
rect -307 -45100 -306 -40970
rect 14 -45100 15 -40970
rect -307 -45101 15 -45100
rect -198 -45499 -94 -45101
rect 282 -45152 302 -40918
rect 366 -45152 386 -40918
rect 282 -45448 386 -45152
rect -307 -45500 15 -45499
rect -307 -49630 -306 -45500
rect 14 -49630 15 -45500
rect -307 -49631 15 -49630
rect -198 -50029 -94 -49631
rect 282 -49682 302 -45448
rect 366 -49682 386 -45448
rect 282 -49978 386 -49682
rect -307 -50030 15 -50029
rect -307 -54160 -306 -50030
rect 14 -54160 15 -50030
rect -307 -54161 15 -54160
rect -198 -54559 -94 -54161
rect 282 -54212 302 -49978
rect 366 -54212 386 -49978
rect 282 -54508 386 -54212
rect -307 -54560 15 -54559
rect -307 -58690 -306 -54560
rect 14 -58690 15 -54560
rect -307 -58691 15 -58690
rect -198 -59089 -94 -58691
rect 282 -58742 302 -54508
rect 366 -58742 386 -54508
rect 282 -59038 386 -58742
rect -307 -59090 15 -59089
rect -307 -63220 -306 -59090
rect 14 -63220 15 -59090
rect -307 -63221 15 -63220
rect -198 -63619 -94 -63221
rect 282 -63272 302 -59038
rect 366 -63272 386 -59038
rect 282 -63568 386 -63272
rect -307 -63620 15 -63619
rect -307 -67750 -306 -63620
rect 14 -67750 15 -63620
rect -307 -67751 15 -67750
rect -198 -68149 -94 -67751
rect 282 -67802 302 -63568
rect 366 -67802 386 -63568
rect 282 -68098 386 -67802
rect -307 -68150 15 -68149
rect -307 -72280 -306 -68150
rect 14 -72280 15 -68150
rect -307 -72281 15 -72280
rect -198 -72679 -94 -72281
rect 282 -72332 302 -68098
rect 366 -72332 386 -68098
rect 282 -72628 386 -72332
rect -307 -72680 15 -72679
rect -307 -76810 -306 -72680
rect 14 -76810 15 -72680
rect -307 -76811 15 -76810
rect -198 -77209 -94 -76811
rect 282 -76862 302 -72628
rect 366 -76862 386 -72628
rect 282 -77158 386 -76862
rect -307 -77210 15 -77209
rect -307 -81340 -306 -77210
rect 14 -81340 15 -77210
rect -307 -81341 15 -81340
rect -198 -81739 -94 -81341
rect 282 -81392 302 -77158
rect 366 -81392 386 -77158
rect 282 -81688 386 -81392
rect -307 -81740 15 -81739
rect -307 -85870 -306 -81740
rect 14 -85870 15 -81740
rect -307 -85871 15 -85870
rect -198 -86269 -94 -85871
rect 282 -85922 302 -81688
rect 366 -85922 386 -81688
rect 282 -86218 386 -85922
rect -307 -86270 15 -86269
rect -307 -90400 -306 -86270
rect 14 -90400 15 -86270
rect -307 -90401 15 -90400
rect -198 -90799 -94 -90401
rect 282 -90452 302 -86218
rect 366 -90452 386 -86218
rect 282 -90748 386 -90452
rect -307 -90800 15 -90799
rect -307 -94930 -306 -90800
rect 14 -94930 15 -90800
rect -307 -94931 15 -94930
rect -198 -95329 -94 -94931
rect 282 -94982 302 -90748
rect 366 -94982 386 -90748
rect 282 -95278 386 -94982
rect -307 -95330 15 -95329
rect -307 -99460 -306 -95330
rect 14 -99460 15 -95330
rect -307 -99461 15 -99460
rect -198 -99859 -94 -99461
rect 282 -99512 302 -95278
rect 366 -99512 386 -95278
rect 282 -99808 386 -99512
rect -307 -99860 15 -99859
rect -307 -103990 -306 -99860
rect 14 -103990 15 -99860
rect -307 -103991 15 -103990
rect -198 -104389 -94 -103991
rect 282 -104042 302 -99808
rect 366 -104042 386 -99808
rect 282 -104338 386 -104042
rect -307 -104390 15 -104389
rect -307 -108520 -306 -104390
rect 14 -108520 15 -104390
rect -307 -108521 15 -108520
rect -198 -108919 -94 -108521
rect 282 -108572 302 -104338
rect 366 -108572 386 -104338
rect 282 -108868 386 -108572
rect -307 -108920 15 -108919
rect -307 -113050 -306 -108920
rect 14 -113050 15 -108920
rect -307 -113051 15 -113050
rect -198 -113449 -94 -113051
rect 282 -113102 302 -108868
rect 366 -113102 386 -108868
rect 282 -113398 386 -113102
rect -307 -113450 15 -113449
rect -307 -117580 -306 -113450
rect 14 -117580 15 -113450
rect -307 -117581 15 -117580
rect -198 -117979 -94 -117581
rect 282 -117632 302 -113398
rect 366 -117632 386 -113398
rect 282 -117928 386 -117632
rect -307 -117980 15 -117979
rect -307 -122110 -306 -117980
rect 14 -122110 15 -117980
rect -307 -122111 15 -122110
rect -198 -122509 -94 -122111
rect 282 -122162 302 -117928
rect 366 -122162 386 -117928
rect 282 -122458 386 -122162
rect -307 -122510 15 -122509
rect -307 -126640 -306 -122510
rect 14 -126640 15 -122510
rect -307 -126641 15 -126640
rect -198 -127039 -94 -126641
rect 282 -126692 302 -122458
rect 366 -126692 386 -122458
rect 282 -126988 386 -126692
rect -307 -127040 15 -127039
rect -307 -131170 -306 -127040
rect 14 -131170 15 -127040
rect -307 -131171 15 -131170
rect -198 -131569 -94 -131171
rect 282 -131222 302 -126988
rect 366 -131222 386 -126988
rect 282 -131518 386 -131222
rect -307 -131570 15 -131569
rect -307 -135700 -306 -131570
rect 14 -135700 15 -131570
rect -307 -135701 15 -135700
rect -198 -136099 -94 -135701
rect 282 -135752 302 -131518
rect 366 -135752 386 -131518
rect 282 -136048 386 -135752
rect -307 -136100 15 -136099
rect -307 -140230 -306 -136100
rect 14 -140230 15 -136100
rect -307 -140231 15 -140230
rect -198 -140629 -94 -140231
rect 282 -140282 302 -136048
rect 366 -140282 386 -136048
rect 282 -140578 386 -140282
rect -307 -140630 15 -140629
rect -307 -144760 -306 -140630
rect 14 -144760 15 -140630
rect -307 -144761 15 -144760
rect -198 -145159 -94 -144761
rect 282 -144812 302 -140578
rect 366 -144812 386 -140578
rect 282 -145108 386 -144812
rect -307 -145160 15 -145159
rect -307 -149290 -306 -145160
rect 14 -149290 15 -145160
rect -307 -149291 15 -149290
rect -198 -149689 -94 -149291
rect 282 -149342 302 -145108
rect 366 -149342 386 -145108
rect 282 -149638 386 -149342
rect -307 -149690 15 -149689
rect -307 -153820 -306 -149690
rect 14 -153820 15 -149690
rect -307 -153821 15 -153820
rect -198 -154219 -94 -153821
rect 282 -153872 302 -149638
rect 366 -153872 386 -149638
rect 282 -154168 386 -153872
rect -307 -154220 15 -154219
rect -307 -158350 -306 -154220
rect 14 -158350 15 -154220
rect -307 -158351 15 -158350
rect -198 -158749 -94 -158351
rect 282 -158402 302 -154168
rect 366 -158402 386 -154168
rect 282 -158698 386 -158402
rect -307 -158750 15 -158749
rect -307 -162880 -306 -158750
rect 14 -162880 15 -158750
rect -307 -162881 15 -162880
rect -198 -163279 -94 -162881
rect 282 -162932 302 -158698
rect 366 -162932 386 -158698
rect 282 -163228 386 -162932
rect -307 -163280 15 -163279
rect -307 -167410 -306 -163280
rect 14 -167410 15 -163280
rect -307 -167411 15 -167410
rect -198 -167809 -94 -167411
rect 282 -167462 302 -163228
rect 366 -167462 386 -163228
rect 282 -167758 386 -167462
rect -307 -167810 15 -167809
rect -307 -171940 -306 -167810
rect 14 -171940 15 -167810
rect -307 -171941 15 -171940
rect -198 -172339 -94 -171941
rect 282 -171992 302 -167758
rect 366 -171992 386 -167758
rect 282 -172288 386 -171992
rect -307 -172340 15 -172339
rect -307 -176470 -306 -172340
rect 14 -176470 15 -172340
rect -307 -176471 15 -176470
rect -198 -176869 -94 -176471
rect 282 -176522 302 -172288
rect 366 -176522 386 -172288
rect 282 -176818 386 -176522
rect -307 -176870 15 -176869
rect -307 -181000 -306 -176870
rect 14 -181000 15 -176870
rect -307 -181001 15 -181000
rect -198 -181399 -94 -181001
rect 282 -181052 302 -176818
rect 366 -181052 386 -176818
rect 282 -181348 386 -181052
rect -307 -181400 15 -181399
rect -307 -185530 -306 -181400
rect 14 -185530 15 -181400
rect -307 -185531 15 -185530
rect -198 -185929 -94 -185531
rect 282 -185582 302 -181348
rect 366 -185582 386 -181348
rect 282 -185878 386 -185582
rect -307 -185930 15 -185929
rect -307 -190060 -306 -185930
rect 14 -190060 15 -185930
rect -307 -190061 15 -190060
rect -198 -190459 -94 -190061
rect 282 -190112 302 -185878
rect 366 -190112 386 -185878
rect 282 -190408 386 -190112
rect -307 -190460 15 -190459
rect -307 -194590 -306 -190460
rect 14 -194590 15 -190460
rect -307 -194591 15 -194590
rect -198 -194989 -94 -194591
rect 282 -194642 302 -190408
rect 366 -194642 386 -190408
rect 282 -194938 386 -194642
rect -307 -194990 15 -194989
rect -307 -199120 -306 -194990
rect 14 -199120 15 -194990
rect -307 -199121 15 -199120
rect -198 -199519 -94 -199121
rect 282 -199172 302 -194938
rect 366 -199172 386 -194938
rect 282 -199468 386 -199172
rect -307 -199520 15 -199519
rect -307 -203650 -306 -199520
rect 14 -203650 15 -199520
rect -307 -203651 15 -203650
rect -198 -204049 -94 -203651
rect 282 -203702 302 -199468
rect 366 -203702 386 -199468
rect 282 -203998 386 -203702
rect -307 -204050 15 -204049
rect -307 -208180 -306 -204050
rect 14 -208180 15 -204050
rect -307 -208181 15 -208180
rect -198 -208579 -94 -208181
rect 282 -208232 302 -203998
rect 366 -208232 386 -203998
rect 282 -208528 386 -208232
rect -307 -208580 15 -208579
rect -307 -212710 -306 -208580
rect 14 -212710 15 -208580
rect -307 -212711 15 -212710
rect -198 -213109 -94 -212711
rect 282 -212762 302 -208528
rect 366 -212762 386 -208528
rect 282 -213058 386 -212762
rect -307 -213110 15 -213109
rect -307 -217240 -306 -213110
rect 14 -217240 15 -213110
rect -307 -217241 15 -217240
rect -198 -217639 -94 -217241
rect 282 -217292 302 -213058
rect 366 -217292 386 -213058
rect 282 -217588 386 -217292
rect -307 -217640 15 -217639
rect -307 -221770 -306 -217640
rect 14 -221770 15 -217640
rect -307 -221771 15 -221770
rect -198 -222169 -94 -221771
rect 282 -221822 302 -217588
rect 366 -221822 386 -217588
rect 282 -222118 386 -221822
rect -307 -222170 15 -222169
rect -307 -226300 -306 -222170
rect 14 -226300 15 -222170
rect -307 -226301 15 -226300
rect -198 -226699 -94 -226301
rect 282 -226352 302 -222118
rect 366 -226352 386 -222118
rect 282 -226648 386 -226352
rect -307 -226700 15 -226699
rect -307 -230830 -306 -226700
rect 14 -230830 15 -226700
rect -307 -230831 15 -230830
rect -198 -231229 -94 -230831
rect 282 -230882 302 -226648
rect 366 -230882 386 -226648
rect 282 -231178 386 -230882
rect -307 -231230 15 -231229
rect -307 -235360 -306 -231230
rect 14 -235360 15 -231230
rect -307 -235361 15 -235360
rect -198 -235759 -94 -235361
rect 282 -235412 302 -231178
rect 366 -235412 386 -231178
rect 282 -235708 386 -235412
rect -307 -235760 15 -235759
rect -307 -239890 -306 -235760
rect 14 -239890 15 -235760
rect -307 -239891 15 -239890
rect -198 -240289 -94 -239891
rect 282 -239942 302 -235708
rect 366 -239942 386 -235708
rect 282 -240238 386 -239942
rect -307 -240290 15 -240289
rect -307 -244420 -306 -240290
rect 14 -244420 15 -240290
rect -307 -244421 15 -244420
rect -198 -244819 -94 -244421
rect 282 -244472 302 -240238
rect 366 -244472 386 -240238
rect 282 -244768 386 -244472
rect -307 -244820 15 -244819
rect -307 -248950 -306 -244820
rect 14 -248950 15 -244820
rect -307 -248951 15 -248950
rect -198 -249349 -94 -248951
rect 282 -249002 302 -244768
rect 366 -249002 386 -244768
rect 282 -249298 386 -249002
rect -307 -249350 15 -249349
rect -307 -253480 -306 -249350
rect 14 -253480 15 -249350
rect -307 -253481 15 -253480
rect -198 -253879 -94 -253481
rect 282 -253532 302 -249298
rect 366 -253532 386 -249298
rect 282 -253828 386 -253532
rect -307 -253880 15 -253879
rect -307 -258010 -306 -253880
rect 14 -258010 15 -253880
rect -307 -258011 15 -258010
rect -198 -258409 -94 -258011
rect 282 -258062 302 -253828
rect 366 -258062 386 -253828
rect 282 -258358 386 -258062
rect -307 -258410 15 -258409
rect -307 -262540 -306 -258410
rect 14 -262540 15 -258410
rect -307 -262541 15 -262540
rect -198 -262939 -94 -262541
rect 282 -262592 302 -258358
rect 366 -262592 386 -258358
rect 282 -262888 386 -262592
rect -307 -262940 15 -262939
rect -307 -267070 -306 -262940
rect 14 -267070 15 -262940
rect -307 -267071 15 -267070
rect -198 -267469 -94 -267071
rect 282 -267122 302 -262888
rect 366 -267122 386 -262888
rect 282 -267418 386 -267122
rect -307 -267470 15 -267469
rect -307 -271600 -306 -267470
rect 14 -271600 15 -267470
rect -307 -271601 15 -271600
rect -198 -271999 -94 -271601
rect 282 -271652 302 -267418
rect 366 -271652 386 -267418
rect 282 -271948 386 -271652
rect -307 -272000 15 -271999
rect -307 -276130 -306 -272000
rect 14 -276130 15 -272000
rect -307 -276131 15 -276130
rect -198 -276529 -94 -276131
rect 282 -276182 302 -271948
rect 366 -276182 386 -271948
rect 282 -276478 386 -276182
rect -307 -276530 15 -276529
rect -307 -280660 -306 -276530
rect 14 -280660 15 -276530
rect -307 -280661 15 -280660
rect -198 -281059 -94 -280661
rect 282 -280712 302 -276478
rect 366 -280712 386 -276478
rect 282 -281008 386 -280712
rect -307 -281060 15 -281059
rect -307 -285190 -306 -281060
rect 14 -285190 15 -281060
rect -307 -285191 15 -285190
rect -198 -285589 -94 -285191
rect 282 -285242 302 -281008
rect 366 -285242 386 -281008
rect 282 -285538 386 -285242
rect -307 -285590 15 -285589
rect -307 -289720 -306 -285590
rect 14 -289720 15 -285590
rect -307 -289721 15 -289720
rect -198 -289920 -94 -289721
rect 282 -289772 302 -285538
rect 366 -289772 386 -285538
rect 282 -289920 386 -289772
<< properties >>
string FIXED_BBOX -386 285510 94 289800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 128 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
