magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -386 17972 386 18000
rect -386 13738 302 17972
rect 366 13738 386 17972
rect -386 13710 386 13738
rect -386 13442 386 13470
rect -386 9208 302 13442
rect 366 9208 386 13442
rect -386 9180 386 9208
rect -386 8912 386 8940
rect -386 4678 302 8912
rect 366 4678 386 8912
rect -386 4650 386 4678
rect -386 4382 386 4410
rect -386 148 302 4382
rect 366 148 386 4382
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -4382 302 -148
rect 366 -4382 386 -148
rect -386 -4410 386 -4382
rect -386 -4678 386 -4650
rect -386 -8912 302 -4678
rect 366 -8912 386 -4678
rect -386 -8940 386 -8912
rect -386 -9208 386 -9180
rect -386 -13442 302 -9208
rect 366 -13442 386 -9208
rect -386 -13470 386 -13442
rect -386 -13738 386 -13710
rect -386 -17972 302 -13738
rect 366 -17972 386 -13738
rect -386 -18000 386 -17972
<< via3 >>
rect 302 13738 366 17972
rect 302 9208 366 13442
rect 302 4678 366 8912
rect 302 148 366 4382
rect 302 -4382 366 -148
rect 302 -8912 366 -4678
rect 302 -13442 366 -9208
rect 302 -17972 366 -13738
<< mimcap >>
rect -346 17920 54 17960
rect -346 13790 -306 17920
rect 14 13790 54 17920
rect -346 13750 54 13790
rect -346 13390 54 13430
rect -346 9260 -306 13390
rect 14 9260 54 13390
rect -346 9220 54 9260
rect -346 8860 54 8900
rect -346 4730 -306 8860
rect 14 4730 54 8860
rect -346 4690 54 4730
rect -346 4330 54 4370
rect -346 200 -306 4330
rect 14 200 54 4330
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -4330 -306 -200
rect 14 -4330 54 -200
rect -346 -4370 54 -4330
rect -346 -4730 54 -4690
rect -346 -8860 -306 -4730
rect 14 -8860 54 -4730
rect -346 -8900 54 -8860
rect -346 -9260 54 -9220
rect -346 -13390 -306 -9260
rect 14 -13390 54 -9260
rect -346 -13430 54 -13390
rect -346 -13790 54 -13750
rect -346 -17920 -306 -13790
rect 14 -17920 54 -13790
rect -346 -17960 54 -17920
<< mimcapcontact >>
rect -306 13790 14 17920
rect -306 9260 14 13390
rect -306 4730 14 8860
rect -306 200 14 4330
rect -306 -4330 14 -200
rect -306 -8860 14 -4730
rect -306 -13390 14 -9260
rect -306 -17920 14 -13790
<< metal4 >>
rect -198 17921 -94 18120
rect 282 17972 386 18120
rect -307 17920 15 17921
rect -307 13790 -306 17920
rect 14 13790 15 17920
rect -307 13789 15 13790
rect -198 13391 -94 13789
rect 282 13738 302 17972
rect 366 13738 386 17972
rect 282 13442 386 13738
rect -307 13390 15 13391
rect -307 9260 -306 13390
rect 14 9260 15 13390
rect -307 9259 15 9260
rect -198 8861 -94 9259
rect 282 9208 302 13442
rect 366 9208 386 13442
rect 282 8912 386 9208
rect -307 8860 15 8861
rect -307 4730 -306 8860
rect 14 4730 15 8860
rect -307 4729 15 4730
rect -198 4331 -94 4729
rect 282 4678 302 8912
rect 366 4678 386 8912
rect 282 4382 386 4678
rect -307 4330 15 4331
rect -307 200 -306 4330
rect 14 200 15 4330
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 4382
rect 366 148 386 4382
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -4330 -306 -200
rect 14 -4330 15 -200
rect -307 -4331 15 -4330
rect -198 -4729 -94 -4331
rect 282 -4382 302 -148
rect 366 -4382 386 -148
rect 282 -4678 386 -4382
rect -307 -4730 15 -4729
rect -307 -8860 -306 -4730
rect 14 -8860 15 -4730
rect -307 -8861 15 -8860
rect -198 -9259 -94 -8861
rect 282 -8912 302 -4678
rect 366 -8912 386 -4678
rect 282 -9208 386 -8912
rect -307 -9260 15 -9259
rect -307 -13390 -306 -9260
rect 14 -13390 15 -9260
rect -307 -13391 15 -13390
rect -198 -13789 -94 -13391
rect 282 -13442 302 -9208
rect 366 -13442 386 -9208
rect 282 -13738 386 -13442
rect -307 -13790 15 -13789
rect -307 -17920 -306 -13790
rect 14 -17920 15 -13790
rect -307 -17921 15 -17920
rect -198 -18120 -94 -17921
rect 282 -17972 302 -13738
rect 366 -17972 386 -13738
rect 282 -18120 386 -17972
<< properties >>
string FIXED_BBOX -386 13710 94 18000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 1 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
