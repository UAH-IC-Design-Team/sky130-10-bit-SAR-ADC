magic
tech sky130A
magscale 1 2
timestamp 1666311401
<< metal4 >>
rect 200 0 300 38000
rect 600 0 700 38000
rect 1200 0 1300 38000
rect 1600 0 1700 38000
rect 2200 0 2300 38000
rect 2600 0 2700 38000
rect 3200 0 3300 38000
rect 3600 0 3700 38000
rect 4200 0 4300 38000
rect 4600 0 4700 38000
rect 5200 0 5300 38000
rect 5600 0 5700 38000
rect 6200 0 6300 38000
rect 6600 0 6700 38000
rect 7200 0 7300 38000
rect 7600 0 7700 38000
rect 8200 0 8300 38000
rect 8600 0 8700 38000
rect 9200 0 9300 38000
rect 9600 0 9700 38000
rect 10200 0 10300 38000
rect 10600 0 10700 38000
rect 11200 0 11300 38000
rect 11600 0 11700 38000
rect 12200 0 12300 38000
rect 12600 0 12700 38000
rect 13200 0 13300 38000
rect 13600 0 13700 38000
rect 14200 0 14300 38000
rect 14600 0 14700 38000
rect 15200 0 15300 38000
rect 15600 0 15700 38000
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  sky130_fd_pr__cap_mim_m3_1_LQSHR5_0
array 0 15 1000 0 7 4800
timestamp 1666311151
transform 1 0 350 0 1 2205
box -350 -2205 349 2205
<< end >>
