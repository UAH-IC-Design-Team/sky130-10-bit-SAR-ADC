magic
tech sky130A
magscale 1 2
timestamp 1665617364
<< error_p >>
rect -50 50 -10 650
rect 10 50 50 650
rect -50 -650 -10 -50
rect 10 -650 50 -50
<< metal3 >>
rect -709 622 -10 650
rect -709 78 -94 622
rect -30 78 -10 622
rect -709 50 -10 78
rect 10 622 709 650
rect 10 78 625 622
rect 689 78 709 622
rect 10 50 709 78
rect -709 -78 -10 -50
rect -709 -622 -94 -78
rect -30 -622 -10 -78
rect -709 -650 -10 -622
rect 10 -78 709 -50
rect 10 -622 625 -78
rect 689 -622 709 -78
rect 10 -650 709 -622
<< via3 >>
rect -94 78 -30 622
rect 625 78 689 622
rect -94 -622 -30 -78
rect 625 -622 689 -78
<< mimcap >>
rect -609 510 -209 550
rect -609 190 -569 510
rect -249 190 -209 510
rect -609 150 -209 190
rect 110 510 510 550
rect 110 190 150 510
rect 470 190 510 510
rect 110 150 510 190
rect -609 -190 -209 -150
rect -609 -510 -569 -190
rect -249 -510 -209 -190
rect -609 -550 -209 -510
rect 110 -190 510 -150
rect 110 -510 150 -190
rect 470 -510 510 -190
rect 110 -550 510 -510
<< mimcapcontact >>
rect -569 190 -249 510
rect 150 190 470 510
rect -569 -510 -249 -190
rect 150 -510 470 -190
<< metal4 >>
rect -461 511 -357 700
rect -141 638 -37 700
rect -141 622 -14 638
rect -570 510 -248 511
rect -570 190 -569 510
rect -249 190 -248 510
rect -570 189 -248 190
rect -461 -189 -357 189
rect -141 78 -94 622
rect -30 78 -14 622
rect 258 511 362 700
rect 578 638 682 700
rect 578 622 705 638
rect 149 510 471 511
rect 149 190 150 510
rect 470 190 471 510
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -510 -569 -190
rect -249 -510 -248 -190
rect -570 -511 -248 -510
rect -461 -700 -357 -511
rect -141 -622 -94 -78
rect -30 -622 -14 -78
rect 258 -189 362 189
rect 578 78 625 622
rect 689 78 705 622
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -510 150 -190
rect 470 -510 471 -190
rect 149 -511 471 -510
rect -141 -638 -14 -622
rect -141 -700 -37 -638
rect 258 -700 362 -511
rect 578 -622 625 -78
rect 689 -622 705 -78
rect 578 -638 705 -622
rect 578 -700 682 -638
<< properties >>
string FIXED_BBOX 10 50 610 650
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
