magic
tech sky130A
magscale 1 2
timestamp 1666649035
<< error_p >>
rect -29 1053 29 1059
rect -29 1019 -17 1053
rect -29 1013 29 1019
rect -29 725 29 731
rect -29 691 -17 725
rect -29 685 29 691
rect -29 617 29 623
rect -29 583 -17 617
rect -29 577 29 583
rect -29 289 29 295
rect -29 255 -17 289
rect -29 249 29 255
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
rect -29 -255 29 -249
rect -29 -289 -17 -255
rect -29 -295 29 -289
rect -29 -583 29 -577
rect -29 -617 -17 -583
rect -29 -623 29 -617
rect -29 -691 29 -685
rect -29 -725 -17 -691
rect -29 -731 29 -725
rect -29 -1019 29 -1013
rect -29 -1053 -17 -1019
rect -29 -1059 29 -1053
<< nwell >>
rect -211 -1191 211 1191
<< pmos >>
rect -15 772 15 972
rect -15 336 15 536
rect -15 -100 15 100
rect -15 -536 15 -336
rect -15 -972 15 -772
<< pdiff >>
rect -73 960 -15 972
rect -73 784 -61 960
rect -27 784 -15 960
rect -73 772 -15 784
rect 15 960 73 972
rect 15 784 27 960
rect 61 784 73 960
rect 15 772 73 784
rect -73 524 -15 536
rect -73 348 -61 524
rect -27 348 -15 524
rect -73 336 -15 348
rect 15 524 73 536
rect 15 348 27 524
rect 61 348 73 524
rect 15 336 73 348
rect -73 88 -15 100
rect -73 -88 -61 88
rect -27 -88 -15 88
rect -73 -100 -15 -88
rect 15 88 73 100
rect 15 -88 27 88
rect 61 -88 73 88
rect 15 -100 73 -88
rect -73 -348 -15 -336
rect -73 -524 -61 -348
rect -27 -524 -15 -348
rect -73 -536 -15 -524
rect 15 -348 73 -336
rect 15 -524 27 -348
rect 61 -524 73 -348
rect 15 -536 73 -524
rect -73 -784 -15 -772
rect -73 -960 -61 -784
rect -27 -960 -15 -784
rect -73 -972 -15 -960
rect 15 -784 73 -772
rect 15 -960 27 -784
rect 61 -960 73 -784
rect 15 -972 73 -960
<< pdiffc >>
rect -61 784 -27 960
rect 27 784 61 960
rect -61 348 -27 524
rect 27 348 61 524
rect -61 -88 -27 88
rect 27 -88 61 88
rect -61 -524 -27 -348
rect 27 -524 61 -348
rect -61 -960 -27 -784
rect 27 -960 61 -784
<< nsubdiff >>
rect -175 1121 -79 1155
rect 79 1121 175 1155
rect -175 1059 -141 1121
rect 141 1059 175 1121
rect -175 -1121 -141 -1059
rect 141 -1121 175 -1059
rect -175 -1155 -79 -1121
rect 79 -1155 175 -1121
<< nsubdiffcont >>
rect -79 1121 79 1155
rect -175 -1059 -141 1059
rect 141 -1059 175 1059
rect -79 -1155 79 -1121
<< poly >>
rect -33 1053 33 1069
rect -33 1019 -17 1053
rect 17 1019 33 1053
rect -33 1003 33 1019
rect -15 972 15 1003
rect -15 741 15 772
rect -33 725 33 741
rect -33 691 -17 725
rect 17 691 33 725
rect -33 675 33 691
rect -33 617 33 633
rect -33 583 -17 617
rect 17 583 33 617
rect -33 567 33 583
rect -15 536 15 567
rect -15 305 15 336
rect -33 289 33 305
rect -33 255 -17 289
rect 17 255 33 289
rect -33 239 33 255
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -15 100 15 131
rect -15 -131 15 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
rect -33 -255 33 -239
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -305 33 -289
rect -15 -336 15 -305
rect -15 -567 15 -536
rect -33 -583 33 -567
rect -33 -617 -17 -583
rect 17 -617 33 -583
rect -33 -633 33 -617
rect -33 -691 33 -675
rect -33 -725 -17 -691
rect 17 -725 33 -691
rect -33 -741 33 -725
rect -15 -772 15 -741
rect -15 -1003 15 -972
rect -33 -1019 33 -1003
rect -33 -1053 -17 -1019
rect 17 -1053 33 -1019
rect -33 -1069 33 -1053
<< polycont >>
rect -17 1019 17 1053
rect -17 691 17 725
rect -17 583 17 617
rect -17 255 17 289
rect -17 147 17 181
rect -17 -181 17 -147
rect -17 -289 17 -255
rect -17 -617 17 -583
rect -17 -725 17 -691
rect -17 -1053 17 -1019
<< locali >>
rect -175 1121 -79 1155
rect 79 1121 175 1155
rect -175 1059 -141 1121
rect 141 1059 175 1121
rect -33 1019 -17 1053
rect 17 1019 33 1053
rect -61 960 -27 976
rect -61 768 -27 784
rect 27 960 61 976
rect 27 768 61 784
rect -33 691 -17 725
rect 17 691 33 725
rect -33 583 -17 617
rect 17 583 33 617
rect -61 524 -27 540
rect -61 332 -27 348
rect 27 524 61 540
rect 27 332 61 348
rect -33 255 -17 289
rect 17 255 33 289
rect -33 147 -17 181
rect 17 147 33 181
rect -61 88 -27 104
rect -61 -104 -27 -88
rect 27 88 61 104
rect 27 -104 61 -88
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -61 -348 -27 -332
rect -61 -540 -27 -524
rect 27 -348 61 -332
rect 27 -540 61 -524
rect -33 -617 -17 -583
rect 17 -617 33 -583
rect -33 -725 -17 -691
rect 17 -725 33 -691
rect -61 -784 -27 -768
rect -61 -976 -27 -960
rect 27 -784 61 -768
rect 27 -976 61 -960
rect -33 -1053 -17 -1019
rect 17 -1053 33 -1019
rect -175 -1121 -141 -1059
rect 141 -1121 175 -1059
rect -175 -1155 -79 -1121
rect 79 -1155 175 -1121
<< viali >>
rect -17 1019 17 1053
rect -61 784 -27 960
rect 27 784 61 960
rect -17 691 17 725
rect -17 583 17 617
rect -61 348 -27 524
rect 27 348 61 524
rect -17 255 17 289
rect -17 147 17 181
rect -61 -88 -27 88
rect 27 -88 61 88
rect -17 -181 17 -147
rect -17 -289 17 -255
rect -61 -524 -27 -348
rect 27 -524 61 -348
rect -17 -617 17 -583
rect -17 -725 17 -691
rect -61 -960 -27 -784
rect 27 -960 61 -784
rect -17 -1053 17 -1019
<< metal1 >>
rect -29 1053 29 1059
rect -29 1019 -17 1053
rect 17 1019 29 1053
rect -29 1013 29 1019
rect -67 960 -21 972
rect -67 784 -61 960
rect -27 784 -21 960
rect -67 772 -21 784
rect 21 960 67 972
rect 21 784 27 960
rect 61 784 67 960
rect 21 772 67 784
rect -29 725 29 731
rect -29 691 -17 725
rect 17 691 29 725
rect -29 685 29 691
rect -29 617 29 623
rect -29 583 -17 617
rect 17 583 29 617
rect -29 577 29 583
rect -67 524 -21 536
rect -67 348 -61 524
rect -27 348 -21 524
rect -67 336 -21 348
rect 21 524 67 536
rect 21 348 27 524
rect 61 348 67 524
rect 21 336 67 348
rect -29 289 29 295
rect -29 255 -17 289
rect 17 255 29 289
rect -29 249 29 255
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -67 88 -21 100
rect -67 -88 -61 88
rect -27 -88 -21 88
rect -67 -100 -21 -88
rect 21 88 67 100
rect 21 -88 27 88
rect 61 -88 67 88
rect 21 -100 67 -88
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
rect -29 -255 29 -249
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -295 29 -289
rect -67 -348 -21 -336
rect -67 -524 -61 -348
rect -27 -524 -21 -348
rect -67 -536 -21 -524
rect 21 -348 67 -336
rect 21 -524 27 -348
rect 61 -524 67 -348
rect 21 -536 67 -524
rect -29 -583 29 -577
rect -29 -617 -17 -583
rect 17 -617 29 -583
rect -29 -623 29 -617
rect -29 -691 29 -685
rect -29 -725 -17 -691
rect 17 -725 29 -691
rect -29 -731 29 -725
rect -67 -784 -21 -772
rect -67 -960 -61 -784
rect -27 -960 -21 -784
rect -67 -972 -21 -960
rect 21 -784 67 -772
rect 21 -960 27 -784
rect 61 -960 67 -784
rect 21 -972 67 -960
rect -29 -1019 29 -1013
rect -29 -1053 -17 -1019
rect 17 -1053 29 -1019
rect -29 -1059 29 -1053
<< properties >>
string FIXED_BBOX -158 -1138 158 1138
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
