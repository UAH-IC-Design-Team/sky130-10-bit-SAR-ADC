magic
tech sky130A
magscale 1 2
timestamp 1666553528
<< nwell >>
rect -451 -265 449 205
<< pmos >>
rect -351 -165 -321 165
rect -255 -165 -225 165
rect -159 -165 -129 165
rect -63 -165 -33 165
rect 33 -165 63 165
rect 129 -165 159 165
rect 225 -165 255 165
rect 321 -165 351 165
<< pdiff >>
rect -413 153 -351 165
rect -413 -153 -401 153
rect -367 -153 -351 153
rect -413 -165 -351 -153
rect -321 153 -255 165
rect -321 -153 -305 153
rect -271 -153 -255 153
rect -321 -165 -255 -153
rect -225 153 -159 165
rect -225 -153 -209 153
rect -175 -153 -159 153
rect -225 -165 -159 -153
rect -129 153 -63 165
rect -129 -153 -113 153
rect -79 -153 -63 153
rect -129 -165 -63 -153
rect -33 153 33 165
rect -33 -153 -17 153
rect 17 -153 33 153
rect -33 -165 33 -153
rect 63 153 129 165
rect 63 -153 79 153
rect 113 -153 129 153
rect 63 -165 129 -153
rect 159 153 225 165
rect 159 -153 175 153
rect 209 -153 225 153
rect 159 -165 225 -153
rect 255 153 321 165
rect 255 -153 271 153
rect 305 -153 321 153
rect 255 -165 321 -153
rect 351 153 413 165
rect 351 -153 367 153
rect 401 -153 413 153
rect 351 -165 413 -153
<< pdiffc >>
rect -401 -153 -367 153
rect -305 -153 -271 153
rect -209 -153 -175 153
rect -113 -153 -79 153
rect -17 -153 17 153
rect 79 -153 113 153
rect 175 -153 209 153
rect 271 -153 305 153
rect 367 -153 401 153
<< poly >>
rect -351 165 -321 191
rect -255 165 -225 195
rect -159 165 -129 191
rect -63 165 -33 195
rect 33 165 63 191
rect 129 165 159 195
rect 225 165 255 191
rect 321 165 351 195
rect -351 -196 -321 -165
rect -255 -196 -225 -165
rect -159 -196 -129 -165
rect -63 -196 -33 -165
rect 33 -196 63 -165
rect 129 -196 159 -165
rect 225 -196 255 -165
rect 321 -196 351 -165
rect -377 -212 383 -196
rect -377 -246 -353 -212
rect -319 -246 -257 -212
rect -223 -246 -161 -212
rect -127 -246 -67 -212
rect -33 -246 31 -212
rect 65 -246 123 -212
rect 157 -246 223 -212
rect 257 -246 313 -212
rect 347 -246 383 -212
rect -377 -262 383 -246
<< polycont >>
rect -353 -246 -319 -212
rect -257 -246 -223 -212
rect -161 -246 -127 -212
rect -67 -246 -33 -212
rect 31 -246 65 -212
rect 123 -246 157 -212
rect 223 -246 257 -212
rect 313 -246 347 -212
<< locali >>
rect -401 153 -367 169
rect -401 -169 -367 -153
rect -305 153 -271 169
rect -305 -169 -271 -153
rect -209 153 -175 169
rect -209 -169 -175 -153
rect -113 153 -79 169
rect -113 -169 -79 -153
rect -17 153 17 169
rect -17 -169 17 -153
rect 79 153 113 169
rect 79 -169 113 -153
rect 175 153 209 169
rect 175 -169 209 -153
rect 271 153 305 169
rect 271 -169 305 -153
rect 367 153 401 169
rect 367 -169 401 -153
rect -377 -246 -353 -212
rect -319 -246 -257 -212
rect -223 -246 -161 -212
rect -127 -246 -67 -212
rect -33 -246 31 -212
rect 65 -246 123 -212
rect 157 -246 223 -212
rect 257 -246 313 -212
rect 347 -246 383 -212
<< viali >>
rect -401 44 -367 136
rect -305 -136 -271 -44
rect -209 44 -175 136
rect -113 -136 -79 -44
rect -17 44 17 136
rect 79 -136 113 -44
rect 175 44 209 136
rect 271 -136 305 -44
rect 367 44 401 136
rect -353 -246 -319 -212
rect -257 -246 -223 -212
rect -161 -246 -127 -212
rect -67 -246 -33 -212
rect 31 -246 65 -212
rect 123 -246 157 -212
rect 223 -246 257 -212
rect 313 -246 347 -212
<< metal1 >>
rect -407 136 -361 148
rect -407 44 -401 136
rect -367 44 -361 136
rect -407 32 -361 44
rect -215 136 -169 148
rect -215 44 -209 136
rect -175 44 -169 136
rect -215 32 -169 44
rect -23 136 23 148
rect -23 44 -17 136
rect 17 44 23 136
rect -23 32 23 44
rect 169 136 215 148
rect 169 44 175 136
rect 209 44 215 136
rect 169 32 215 44
rect 361 136 407 148
rect 361 44 367 136
rect 401 44 407 136
rect 361 32 407 44
rect -311 -44 -265 -32
rect -311 -136 -305 -44
rect -271 -136 -265 -44
rect -311 -148 -265 -136
rect -119 -44 -73 -32
rect -119 -136 -113 -44
rect -79 -136 -73 -44
rect -119 -148 -73 -136
rect 73 -44 119 -32
rect 73 -136 79 -44
rect 113 -136 119 -44
rect 73 -148 119 -136
rect 265 -44 311 -32
rect 265 -136 271 -44
rect 305 -136 311 -44
rect 265 -148 311 -136
rect -377 -212 383 -206
rect -377 -246 -353 -212
rect -319 -246 -257 -212
rect -223 -246 -161 -212
rect -127 -246 -67 -212
rect -33 -246 31 -212
rect 65 -246 123 -212
rect 157 -246 223 -212
rect 257 -246 313 -212
rect 347 -246 383 -212
rect -377 -252 383 -246
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
