magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< error_p >>
rect -70 13580 -10 17990
rect 10 13580 70 17990
rect -70 9070 -10 13480
rect 10 9070 70 13480
rect -70 4560 -10 8970
rect 10 4560 70 8970
rect -70 50 -10 4460
rect 10 50 70 4460
rect -70 -4460 -10 -50
rect 10 -4460 70 -50
rect -70 -8970 -10 -4560
rect 10 -8970 70 -4560
rect -70 -13480 -10 -9070
rect 10 -13480 70 -9070
rect -70 -17990 -10 -13580
rect 10 -17990 70 -13580
<< metal3 >>
rect -709 17962 -10 17990
rect -709 13608 -94 17962
rect -30 13608 -10 17962
rect -709 13580 -10 13608
rect 10 17962 709 17990
rect 10 13608 625 17962
rect 689 13608 709 17962
rect 10 13580 709 13608
rect -709 13452 -10 13480
rect -709 9098 -94 13452
rect -30 9098 -10 13452
rect -709 9070 -10 9098
rect 10 13452 709 13480
rect 10 9098 625 13452
rect 689 9098 709 13452
rect 10 9070 709 9098
rect -709 8942 -10 8970
rect -709 4588 -94 8942
rect -30 4588 -10 8942
rect -709 4560 -10 4588
rect 10 8942 709 8970
rect 10 4588 625 8942
rect 689 4588 709 8942
rect 10 4560 709 4588
rect -709 4432 -10 4460
rect -709 78 -94 4432
rect -30 78 -10 4432
rect -709 50 -10 78
rect 10 4432 709 4460
rect 10 78 625 4432
rect 689 78 709 4432
rect 10 50 709 78
rect -709 -78 -10 -50
rect -709 -4432 -94 -78
rect -30 -4432 -10 -78
rect -709 -4460 -10 -4432
rect 10 -78 709 -50
rect 10 -4432 625 -78
rect 689 -4432 709 -78
rect 10 -4460 709 -4432
rect -709 -4588 -10 -4560
rect -709 -8942 -94 -4588
rect -30 -8942 -10 -4588
rect -709 -8970 -10 -8942
rect 10 -4588 709 -4560
rect 10 -8942 625 -4588
rect 689 -8942 709 -4588
rect 10 -8970 709 -8942
rect -709 -9098 -10 -9070
rect -709 -13452 -94 -9098
rect -30 -13452 -10 -9098
rect -709 -13480 -10 -13452
rect 10 -9098 709 -9070
rect 10 -13452 625 -9098
rect 689 -13452 709 -9098
rect 10 -13480 709 -13452
rect -709 -13608 -10 -13580
rect -709 -17962 -94 -13608
rect -30 -17962 -10 -13608
rect -709 -17990 -10 -17962
rect 10 -13608 709 -13580
rect 10 -17962 625 -13608
rect 689 -17962 709 -13608
rect 10 -17990 709 -17962
<< via3 >>
rect -94 13608 -30 17962
rect 625 13608 689 17962
rect -94 9098 -30 13452
rect 625 9098 689 13452
rect -94 4588 -30 8942
rect 625 4588 689 8942
rect -94 78 -30 4432
rect 625 78 689 4432
rect -94 -4432 -30 -78
rect 625 -4432 689 -78
rect -94 -8942 -30 -4588
rect 625 -8942 689 -4588
rect -94 -13452 -30 -9098
rect 625 -13452 689 -9098
rect -94 -17962 -30 -13608
rect 625 -17962 689 -13608
<< mimcap >>
rect -609 17850 -209 17890
rect -609 13720 -569 17850
rect -249 13720 -209 17850
rect -609 13680 -209 13720
rect 110 17850 510 17890
rect 110 13720 150 17850
rect 470 13720 510 17850
rect 110 13680 510 13720
rect -609 13340 -209 13380
rect -609 9210 -569 13340
rect -249 9210 -209 13340
rect -609 9170 -209 9210
rect 110 13340 510 13380
rect 110 9210 150 13340
rect 470 9210 510 13340
rect 110 9170 510 9210
rect -609 8830 -209 8870
rect -609 4700 -569 8830
rect -249 4700 -209 8830
rect -609 4660 -209 4700
rect 110 8830 510 8870
rect 110 4700 150 8830
rect 470 4700 510 8830
rect 110 4660 510 4700
rect -609 4320 -209 4360
rect -609 190 -569 4320
rect -249 190 -209 4320
rect -609 150 -209 190
rect 110 4320 510 4360
rect 110 190 150 4320
rect 470 190 510 4320
rect 110 150 510 190
rect -609 -190 -209 -150
rect -609 -4320 -569 -190
rect -249 -4320 -209 -190
rect -609 -4360 -209 -4320
rect 110 -190 510 -150
rect 110 -4320 150 -190
rect 470 -4320 510 -190
rect 110 -4360 510 -4320
rect -609 -4700 -209 -4660
rect -609 -8830 -569 -4700
rect -249 -8830 -209 -4700
rect -609 -8870 -209 -8830
rect 110 -4700 510 -4660
rect 110 -8830 150 -4700
rect 470 -8830 510 -4700
rect 110 -8870 510 -8830
rect -609 -9210 -209 -9170
rect -609 -13340 -569 -9210
rect -249 -13340 -209 -9210
rect -609 -13380 -209 -13340
rect 110 -9210 510 -9170
rect 110 -13340 150 -9210
rect 470 -13340 510 -9210
rect 110 -13380 510 -13340
rect -609 -13720 -209 -13680
rect -609 -17850 -569 -13720
rect -249 -17850 -209 -13720
rect -609 -17890 -209 -17850
rect 110 -13720 510 -13680
rect 110 -17850 150 -13720
rect 470 -17850 510 -13720
rect 110 -17890 510 -17850
<< mimcapcontact >>
rect -569 13720 -249 17850
rect 150 13720 470 17850
rect -569 9210 -249 13340
rect 150 9210 470 13340
rect -569 4700 -249 8830
rect 150 4700 470 8830
rect -569 190 -249 4320
rect 150 190 470 4320
rect -569 -4320 -249 -190
rect 150 -4320 470 -190
rect -569 -8830 -249 -4700
rect 150 -8830 470 -4700
rect -569 -13340 -249 -9210
rect 150 -13340 470 -9210
rect -569 -17850 -249 -13720
rect 150 -17850 470 -13720
<< metal4 >>
rect -461 17851 -357 18040
rect -141 17978 -37 18040
rect -141 17962 -14 17978
rect -570 17850 -248 17851
rect -570 13720 -569 17850
rect -249 13720 -248 17850
rect -570 13719 -248 13720
rect -461 13341 -357 13719
rect -141 13608 -94 17962
rect -30 13608 -14 17962
rect 258 17851 362 18040
rect 578 17978 682 18040
rect 578 17962 705 17978
rect 149 17850 471 17851
rect 149 13720 150 17850
rect 470 13720 471 17850
rect 149 13719 471 13720
rect -141 13592 -14 13608
rect -141 13468 -37 13592
rect -141 13452 -14 13468
rect -570 13340 -248 13341
rect -570 9210 -569 13340
rect -249 9210 -248 13340
rect -570 9209 -248 9210
rect -461 8831 -357 9209
rect -141 9098 -94 13452
rect -30 9098 -14 13452
rect 258 13341 362 13719
rect 578 13608 625 17962
rect 689 13608 705 17962
rect 578 13592 705 13608
rect 578 13468 682 13592
rect 578 13452 705 13468
rect 149 13340 471 13341
rect 149 9210 150 13340
rect 470 9210 471 13340
rect 149 9209 471 9210
rect -141 9082 -14 9098
rect -141 8958 -37 9082
rect -141 8942 -14 8958
rect -570 8830 -248 8831
rect -570 4700 -569 8830
rect -249 4700 -248 8830
rect -570 4699 -248 4700
rect -461 4321 -357 4699
rect -141 4588 -94 8942
rect -30 4588 -14 8942
rect 258 8831 362 9209
rect 578 9098 625 13452
rect 689 9098 705 13452
rect 578 9082 705 9098
rect 578 8958 682 9082
rect 578 8942 705 8958
rect 149 8830 471 8831
rect 149 4700 150 8830
rect 470 4700 471 8830
rect 149 4699 471 4700
rect -141 4572 -14 4588
rect -141 4448 -37 4572
rect -141 4432 -14 4448
rect -570 4320 -248 4321
rect -570 190 -569 4320
rect -249 190 -248 4320
rect -570 189 -248 190
rect -461 -189 -357 189
rect -141 78 -94 4432
rect -30 78 -14 4432
rect 258 4321 362 4699
rect 578 4588 625 8942
rect 689 4588 705 8942
rect 578 4572 705 4588
rect 578 4448 682 4572
rect 578 4432 705 4448
rect 149 4320 471 4321
rect 149 190 150 4320
rect 470 190 471 4320
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -4320 -569 -190
rect -249 -4320 -248 -190
rect -570 -4321 -248 -4320
rect -461 -4699 -357 -4321
rect -141 -4432 -94 -78
rect -30 -4432 -14 -78
rect 258 -189 362 189
rect 578 78 625 4432
rect 689 78 705 4432
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -4320 150 -190
rect 470 -4320 471 -190
rect 149 -4321 471 -4320
rect -141 -4448 -14 -4432
rect -141 -4572 -37 -4448
rect -141 -4588 -14 -4572
rect -570 -4700 -248 -4699
rect -570 -8830 -569 -4700
rect -249 -8830 -248 -4700
rect -570 -8831 -248 -8830
rect -461 -9209 -357 -8831
rect -141 -8942 -94 -4588
rect -30 -8942 -14 -4588
rect 258 -4699 362 -4321
rect 578 -4432 625 -78
rect 689 -4432 705 -78
rect 578 -4448 705 -4432
rect 578 -4572 682 -4448
rect 578 -4588 705 -4572
rect 149 -4700 471 -4699
rect 149 -8830 150 -4700
rect 470 -8830 471 -4700
rect 149 -8831 471 -8830
rect -141 -8958 -14 -8942
rect -141 -9082 -37 -8958
rect -141 -9098 -14 -9082
rect -570 -9210 -248 -9209
rect -570 -13340 -569 -9210
rect -249 -13340 -248 -9210
rect -570 -13341 -248 -13340
rect -461 -13719 -357 -13341
rect -141 -13452 -94 -9098
rect -30 -13452 -14 -9098
rect 258 -9209 362 -8831
rect 578 -8942 625 -4588
rect 689 -8942 705 -4588
rect 578 -8958 705 -8942
rect 578 -9082 682 -8958
rect 578 -9098 705 -9082
rect 149 -9210 471 -9209
rect 149 -13340 150 -9210
rect 470 -13340 471 -9210
rect 149 -13341 471 -13340
rect -141 -13468 -14 -13452
rect -141 -13592 -37 -13468
rect -141 -13608 -14 -13592
rect -570 -13720 -248 -13719
rect -570 -17850 -569 -13720
rect -249 -17850 -248 -13720
rect -570 -17851 -248 -17850
rect -461 -18040 -357 -17851
rect -141 -17962 -94 -13608
rect -30 -17962 -14 -13608
rect 258 -13719 362 -13341
rect 578 -13452 625 -9098
rect 689 -13452 705 -9098
rect 578 -13468 705 -13452
rect 578 -13592 682 -13468
rect 578 -13608 705 -13592
rect 149 -13720 471 -13719
rect 149 -17850 150 -13720
rect 470 -17850 471 -13720
rect 149 -17851 471 -17850
rect -141 -17978 -14 -17962
rect -141 -18040 -37 -17978
rect 258 -18040 362 -17851
rect 578 -17962 625 -13608
rect 689 -17962 705 -13608
rect 578 -17978 705 -17962
rect 578 -18040 682 -17978
<< properties >>
string FIXED_BBOX 10 13580 610 17990
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 2 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
