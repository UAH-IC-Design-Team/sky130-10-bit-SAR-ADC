magic
tech sky130A
magscale 1 2
timestamp 1668103091
<< nwell >>
rect 65829 66530 66130 66750
rect 65829 66490 66220 66530
rect 67069 66490 67370 66750
rect 68309 66490 68610 66750
rect 69549 66490 69850 66750
rect 70960 66490 71100 66630
rect 64890 63800 65211 66490
rect 65809 63800 66451 66490
rect 67049 63800 67691 66490
rect 68289 63800 68931 66490
rect 69529 63800 70171 66490
rect 70769 66430 71100 66490
rect 70769 63800 71090 66430
rect 65829 63760 66220 63800
rect 65829 63540 66130 63760
rect 67069 63540 67370 63800
rect 68309 63540 68610 63800
rect 69549 63540 69850 63800
rect 65829 39640 66130 39860
rect 65829 39600 66220 39640
rect 67069 39600 67370 39860
rect 68309 39600 68610 39860
rect 69549 39600 69850 39860
rect 64890 36910 65211 39600
rect 65809 36910 66451 39600
rect 67049 36910 67691 39600
rect 68289 36910 68931 39600
rect 69529 36910 70171 39600
rect 70769 36970 71090 39600
rect 70769 36910 71100 36970
rect 65829 36870 66220 36910
rect 65829 36650 66130 36870
rect 67069 36650 67370 36910
rect 68309 36650 68610 36910
rect 69549 36650 69850 36910
rect 70960 36770 71100 36910
<< locali >>
rect 65149 66450 65325 66453
rect 65149 66402 65160 66450
rect 65320 66402 65325 66450
rect 65695 66450 65871 66453
rect 65695 66402 65700 66450
rect 65860 66402 65871 66450
rect 66389 66450 66565 66453
rect 66389 66402 66390 66450
rect 66560 66402 66565 66450
rect 66935 66450 67111 66453
rect 66935 66402 66940 66450
rect 67100 66402 67111 66450
rect 67629 66450 67805 66453
rect 67629 66402 67630 66450
rect 67800 66402 67805 66450
rect 68175 66450 68351 66453
rect 68175 66402 68180 66450
rect 68350 66402 68351 66450
rect 68869 66450 69045 66453
rect 68869 66402 68880 66450
rect 69040 66402 69045 66450
rect 69415 66450 69591 66453
rect 69415 66402 69420 66450
rect 69580 66402 69591 66450
rect 70109 66450 70285 66453
rect 70109 66402 70120 66450
rect 70280 66402 70285 66450
rect 70655 66450 70831 66453
rect 70655 66402 70660 66450
rect 70820 66402 70831 66450
rect 65217 63996 65223 64066
rect 65217 63980 65257 63996
rect 65797 63996 65803 64066
rect 65763 63980 65803 63996
rect 66457 63996 66463 64066
rect 66457 63980 66497 63996
rect 67037 63996 67043 64066
rect 67003 63980 67043 63996
rect 67697 63996 67703 64066
rect 67697 63980 67737 63996
rect 68277 63996 68283 64066
rect 68243 63980 68283 63996
rect 68937 63996 68943 64066
rect 68937 63980 68977 63996
rect 69517 63996 69523 64066
rect 69483 63980 69523 63996
rect 70177 63996 70183 64066
rect 70177 63980 70217 63996
rect 70757 63996 70763 64066
rect 70723 63980 70763 63996
rect 65217 39404 65257 39420
rect 65217 39334 65223 39404
rect 65763 39404 65803 39420
rect 65797 39334 65803 39404
rect 66457 39404 66497 39420
rect 66457 39334 66463 39404
rect 67003 39404 67043 39420
rect 67037 39334 67043 39404
rect 67697 39404 67737 39420
rect 67697 39334 67703 39404
rect 68243 39404 68283 39420
rect 68277 39334 68283 39404
rect 68937 39404 68977 39420
rect 68937 39334 68943 39404
rect 69483 39404 69523 39420
rect 69517 39334 69523 39404
rect 70177 39404 70217 39420
rect 70177 39334 70183 39404
rect 70723 39404 70763 39420
rect 70757 39334 70763 39404
rect 65149 36950 65160 36998
rect 65320 36950 65325 36998
rect 65149 36947 65325 36950
rect 65695 36950 65700 36998
rect 65860 36950 65871 36998
rect 65695 36947 65871 36950
rect 66389 36950 66390 36998
rect 66560 36950 66565 36998
rect 66389 36947 66565 36950
rect 66935 36950 66940 36998
rect 67100 36950 67111 36998
rect 66935 36947 67111 36950
rect 67629 36950 67630 36998
rect 67800 36950 67805 36998
rect 67629 36947 67805 36950
rect 68175 36950 68180 36998
rect 68175 36947 68340 36950
rect 68869 36950 68880 36998
rect 69020 36950 69025 36998
rect 68869 36947 69025 36950
rect 69415 36950 69420 36998
rect 69580 36950 69591 36998
rect 69415 36947 69591 36950
rect 70109 36950 70120 36998
rect 70280 36950 70285 36998
rect 70109 36947 70285 36950
rect 70655 36950 70660 36998
rect 70820 36950 70831 36998
rect 70655 36947 70831 36950
<< viali >>
rect 65210 66550 65270 66690
rect 65750 66550 65810 66680
rect 66450 66550 66510 66680
rect 66990 66550 67050 66680
rect 67690 66560 67750 66680
rect 68230 66570 68290 66690
rect 68930 66560 68990 66680
rect 69470 66560 69530 66680
rect 70170 66560 70230 66680
rect 70710 66560 70770 66680
rect 65160 66370 65320 66450
rect 65700 66370 65860 66450
rect 66390 66370 66560 66450
rect 66940 66370 67100 66450
rect 67630 66370 67800 66450
rect 68180 66370 68350 66450
rect 68880 66370 69040 66450
rect 69420 66370 69580 66450
rect 70120 66370 70280 66450
rect 70660 66370 70820 66450
rect 65223 63996 65257 64110
rect 65763 63996 65797 64110
rect 66463 63996 66497 64110
rect 67003 63996 67037 64110
rect 67703 63996 67737 64110
rect 68243 63996 68277 64110
rect 68943 63996 68977 64110
rect 69483 63996 69517 64110
rect 70183 63996 70217 64110
rect 70723 63996 70757 64110
rect 65210 63600 65270 63740
rect 65750 63610 65810 63740
rect 66450 63610 66510 63740
rect 66990 63610 67050 63740
rect 67690 63610 67750 63730
rect 68230 63600 68290 63720
rect 68930 63610 68990 63730
rect 69470 63610 69530 63730
rect 70170 63610 70230 63730
rect 70710 63610 70770 63730
rect 65210 39660 65270 39800
rect 65750 39660 65810 39790
rect 66450 39660 66510 39790
rect 66990 39660 67050 39790
rect 67690 39670 67750 39790
rect 68230 39680 68290 39800
rect 68930 39670 68990 39790
rect 69470 39670 69530 39790
rect 70170 39670 70230 39790
rect 70710 39670 70770 39790
rect 65223 39290 65257 39404
rect 65763 39290 65797 39404
rect 66463 39290 66497 39404
rect 67003 39290 67037 39404
rect 67703 39290 67737 39404
rect 68243 39290 68277 39404
rect 68943 39290 68977 39404
rect 69483 39290 69517 39404
rect 70183 39290 70217 39404
rect 70723 39290 70757 39404
rect 65160 36950 65320 37030
rect 65700 36950 65860 37030
rect 66390 36950 66560 37030
rect 66940 36950 67100 37030
rect 67630 36950 67800 37030
rect 68180 36950 68340 37030
rect 68880 36950 69020 37030
rect 69420 36950 69580 37030
rect 70120 36950 70280 37030
rect 70660 36950 70820 37030
rect 65210 36710 65270 36850
rect 65750 36720 65810 36850
rect 66450 36720 66510 36850
rect 66990 36720 67050 36850
rect 67690 36720 67750 36840
rect 68230 36710 68290 36830
rect 68930 36720 68990 36840
rect 69470 36720 69530 36840
rect 70170 36720 70230 36840
rect 70710 36720 70770 36840
<< metal1 >>
rect -12200 69340 70770 69400
rect -12200 68340 -12140 69340
rect 600 69240 70230 69300
rect 600 68360 660 69240
rect 26100 69140 69530 69200
rect 26100 68340 26160 69140
rect 38900 69040 68990 69100
rect 38900 68340 38960 69040
rect 46180 68940 68290 69000
rect 46180 68340 46240 68940
rect 49520 68840 67740 68900
rect 49520 68340 49580 68840
rect 51900 68740 67050 68800
rect -13400 67780 -13060 67800
rect -13400 67420 -13380 67780
rect -13220 67420 -13060 67780
rect -13400 67280 -13060 67420
rect -600 67780 -260 67800
rect -600 67420 -580 67780
rect -420 67420 -260 67780
rect -600 67220 -260 67420
rect 24800 67780 25240 67800
rect 24800 67420 24820 67780
rect 24980 67420 25240 67780
rect 24800 67220 25240 67420
rect 37600 67780 38040 67800
rect 37600 67420 37620 67780
rect 37780 67420 38040 67780
rect 37600 67220 38040 67420
rect 46720 67780 47000 67800
rect 46720 67420 46820 67780
rect 46980 67420 47000 67780
rect 46720 67220 47000 67420
rect 50080 67780 50400 67800
rect 50080 67420 50220 67780
rect 50380 67420 50400 67780
rect 51900 67440 51960 68740
rect 57360 68640 66500 68700
rect 57360 68340 57420 68640
rect 60720 68540 65810 68600
rect 60720 68340 60780 68540
rect 63100 68440 65270 68500
rect 57920 67780 58200 67800
rect 50080 67220 50400 67420
rect 57920 67420 58020 67780
rect 58180 67420 58200 67780
rect 52080 67380 52400 67400
rect 52080 67020 52220 67380
rect 52380 67020 52400 67380
rect 57920 67220 58200 67420
rect 61280 67780 61600 67800
rect 61280 67420 61420 67780
rect 61580 67420 61600 67780
rect 63100 67440 63160 68440
rect 61280 67220 61600 67420
rect 63300 67380 63600 67400
rect 52080 67000 52400 67020
rect 63300 67020 63420 67380
rect 63580 67020 63600 67380
rect 63300 67000 63600 67020
rect 65210 66750 65270 68440
rect 65750 66750 65810 68540
rect 66440 66750 66500 68640
rect 66990 66750 67050 68740
rect 67680 66750 67740 68840
rect 68230 66750 68290 68940
rect 68930 66750 68990 69040
rect 69470 66750 69530 69140
rect 70170 66750 70230 69240
rect 70710 66750 70770 69340
rect 580 66400 1220 66460
rect 1400 66400 2060 66460
rect 2240 66400 2280 66460
rect 580 66380 2280 66400
rect 65200 66690 65280 66750
rect 65200 66550 65210 66690
rect 65270 66550 65280 66690
rect 64880 66430 64980 66540
rect 65200 66500 65280 66550
rect 65740 66680 65820 66750
rect 65740 66550 65750 66680
rect 65810 66550 65820 66680
rect 65140 66450 65340 66500
rect 65140 66370 65160 66450
rect 65320 66370 65340 66450
rect 65400 66430 65600 66530
rect 65740 66480 65820 66550
rect 66440 66680 66520 66750
rect 66440 66550 66450 66680
rect 66510 66550 66520 66680
rect 65690 66450 65880 66480
rect 65140 66360 65340 66370
rect 65690 66370 65700 66450
rect 65860 66370 65880 66450
rect 66020 66430 66220 66530
rect 66440 66470 66520 66550
rect 66980 66680 67060 66750
rect 66980 66550 66990 66680
rect 67050 66550 67060 66680
rect 66380 66450 66570 66470
rect 65690 66350 65880 66370
rect 66380 66370 66390 66450
rect 66560 66370 66570 66450
rect 66640 66430 66840 66530
rect 66980 66470 67060 66550
rect 67680 66680 67760 66750
rect 67680 66560 67690 66680
rect 67750 66560 67760 66680
rect 66930 66450 67120 66470
rect 66380 66350 66570 66370
rect 66930 66370 66940 66450
rect 67100 66370 67120 66450
rect 67260 66430 67460 66530
rect 67680 66470 67760 66560
rect 68220 66690 68300 66750
rect 68220 66570 68230 66690
rect 68290 66570 68300 66690
rect 67610 66450 67820 66470
rect 66930 66350 67120 66370
rect 67610 66370 67630 66450
rect 67800 66370 67820 66450
rect 67880 66430 68080 66530
rect 68220 66470 68300 66570
rect 68920 66680 69000 66750
rect 68920 66560 68930 66680
rect 68990 66560 69000 66680
rect 68160 66450 68360 66470
rect 67610 66340 67820 66370
rect 68160 66370 68180 66450
rect 68350 66370 68360 66450
rect 68500 66430 68700 66530
rect 68920 66470 69000 66560
rect 69460 66680 69540 66750
rect 69460 66560 69470 66680
rect 69530 66560 69540 66680
rect 68860 66450 69060 66470
rect 68160 66350 68360 66370
rect 68860 66370 68880 66450
rect 69040 66370 69060 66450
rect 69120 66430 69320 66530
rect 69460 66470 69540 66560
rect 70160 66680 70240 66750
rect 70160 66560 70170 66680
rect 70230 66560 70240 66680
rect 69400 66450 69600 66470
rect 68860 66350 69060 66370
rect 69400 66370 69420 66450
rect 69580 66370 69600 66450
rect 69740 66430 69940 66530
rect 70160 66470 70240 66560
rect 70700 66680 70780 66750
rect 70700 66560 70710 66680
rect 70770 66560 70780 66680
rect 70100 66450 70300 66470
rect 69400 66350 69600 66370
rect 70100 66370 70120 66450
rect 70280 66370 70300 66450
rect 70360 66430 70560 66530
rect 70700 66470 70780 66560
rect 70640 66450 70840 66470
rect 70100 66350 70300 66370
rect 70640 66370 70660 66450
rect 70820 66370 70840 66450
rect 71000 66430 71100 66530
rect 70640 66350 70840 66370
rect 65200 64110 65280 64140
rect 64880 63940 64980 64060
rect 65200 63996 65223 64110
rect 65257 63996 65280 64110
rect 65740 64110 65820 64140
rect 64880 63750 64980 63860
rect 65200 63740 65280 63996
rect 65400 63940 65600 64060
rect 65740 63996 65763 64110
rect 65797 63996 65820 64110
rect 66440 64110 66520 64140
rect 65400 63760 65600 63860
rect 65200 63600 65210 63740
rect 65270 63600 65280 63740
rect 65200 63580 65280 63600
rect 65740 63740 65820 63996
rect 66020 63940 66220 64040
rect 66440 63996 66463 64110
rect 66497 63996 66520 64110
rect 66980 64110 67060 64140
rect 66020 63760 66220 63860
rect 65740 63610 65750 63740
rect 65810 63610 65820 63740
rect 65740 63580 65820 63610
rect 66440 63740 66520 63996
rect 66640 63940 66840 64040
rect 66980 63996 67003 64110
rect 67037 63996 67060 64110
rect 67680 64110 67760 64140
rect 66640 63760 66840 63860
rect 66440 63610 66450 63740
rect 66510 63610 66520 63740
rect 66440 63580 66520 63610
rect 66980 63740 67060 63996
rect 67260 63940 67460 64040
rect 67680 63996 67703 64110
rect 67737 63996 67760 64110
rect 68220 64110 68300 64140
rect 67260 63760 67460 63860
rect 66980 63610 66990 63740
rect 67050 63610 67060 63740
rect 66980 63580 67060 63610
rect 67680 63730 67760 63996
rect 67880 63940 68080 64040
rect 68220 63996 68243 64110
rect 68277 63996 68300 64110
rect 68920 64110 69000 64140
rect 67880 63760 68080 63860
rect 67680 63610 67690 63730
rect 67750 63610 67760 63730
rect 67680 63580 67760 63610
rect 68220 63720 68300 63996
rect 68500 63940 68700 64040
rect 68920 63996 68943 64110
rect 68977 63996 69000 64110
rect 69460 64110 69540 64140
rect 68500 63760 68700 63860
rect 68220 63600 68230 63720
rect 68290 63600 68300 63720
rect 68220 63580 68300 63600
rect 68920 63730 69000 63996
rect 69120 63940 69320 64040
rect 69460 63996 69483 64110
rect 69517 63996 69540 64110
rect 70160 64110 70240 64140
rect 69120 63760 69320 63860
rect 68920 63610 68930 63730
rect 68990 63610 69000 63730
rect 68920 63580 69000 63610
rect 69460 63730 69540 63996
rect 69740 63940 69940 64040
rect 70160 63996 70183 64110
rect 70217 63996 70240 64110
rect 70700 64110 70780 64140
rect 69740 63760 69940 63860
rect 69460 63610 69470 63730
rect 69530 63610 69540 63730
rect 69460 63580 69540 63610
rect 70160 63730 70240 63996
rect 70360 63940 70560 64040
rect 70700 63996 70723 64110
rect 70757 63996 70780 64110
rect 70360 63760 70560 63860
rect 70160 63610 70170 63730
rect 70230 63610 70240 63730
rect 70160 63580 70240 63610
rect 70700 63730 70780 63996
rect 71000 63940 71100 64040
rect 71000 63760 71100 63860
rect 70700 63610 70710 63730
rect 70770 63610 70780 63730
rect 70700 63580 70780 63610
rect 65200 57360 65260 63580
rect 65740 57460 65800 63580
rect 66440 57560 66500 63580
rect 66980 57660 67040 63580
rect 67680 57760 67740 63580
rect 68220 57860 68280 63580
rect 68920 57960 68980 63580
rect 69460 58060 69520 63580
rect 70160 58160 70220 63580
rect 70700 58260 70760 63580
rect 70700 58200 87900 58260
rect 70160 58100 87900 58160
rect 69460 58000 87900 58060
rect 68920 57900 87900 57960
rect 68220 57800 87900 57860
rect 67680 57700 87900 57760
rect 66980 57600 87900 57660
rect 66440 57500 87900 57560
rect 65740 57400 87900 57460
rect 65200 57300 87900 57360
rect 68900 57200 87900 57260
rect 68900 56260 68960 57200
rect 71900 57100 87900 57160
rect 71900 56200 71960 57100
rect 74400 57000 87900 57060
rect 74400 56200 74460 57000
rect 80220 56900 87900 56960
rect 80220 56240 80280 56900
rect 83120 56800 87900 56860
rect 83120 56200 83180 56800
rect 85620 56700 87900 56760
rect 85620 56200 85680 56700
rect 87240 56600 87900 56660
rect 87240 56220 87300 56600
rect 69100 56080 69400 56100
rect 69100 55820 69220 56080
rect 69380 55820 69400 56080
rect 69100 55800 69400 55820
rect 72160 56080 72400 56100
rect 72160 55820 72220 56080
rect 72380 55820 72400 56080
rect 72160 55800 72400 55820
rect 74660 56080 74900 56100
rect 74660 55820 74720 56080
rect 74880 55820 74900 56080
rect 74660 55800 74900 55820
rect 80420 56080 80700 56100
rect 80420 55820 80520 56080
rect 80680 55820 80700 56080
rect 80420 55800 80700 55820
rect 83360 56080 83600 56100
rect 83360 55820 83420 56080
rect 83580 55820 83600 56080
rect 83360 55800 83600 55820
rect 85880 56080 86100 56100
rect 85880 55820 85920 56080
rect 86080 55820 86100 56080
rect 85880 55800 86100 55820
rect 87480 56080 87700 56100
rect 87480 55820 87520 56080
rect 87680 55820 87700 56080
rect 87480 55800 87700 55820
rect 72180 47780 72400 47800
rect 69100 47680 69400 47700
rect 69100 47320 69220 47680
rect 69380 47320 69400 47680
rect 72180 47420 72220 47780
rect 72380 47420 72400 47780
rect 72180 47400 72400 47420
rect 74620 47780 74900 47800
rect 74620 47420 74720 47780
rect 74880 47420 74900 47780
rect 83360 47780 83600 47800
rect 74620 47400 74900 47420
rect 80400 47680 80800 47700
rect 69100 47300 69400 47320
rect 80400 47320 80620 47680
rect 80780 47320 80800 47680
rect 83360 47420 83420 47780
rect 83580 47420 83600 47780
rect 83360 47400 83600 47420
rect 85880 47780 86200 47800
rect 85880 47420 86020 47780
rect 86180 47420 86200 47780
rect 85880 47400 86200 47420
rect 87460 47780 87800 47800
rect 87460 47420 87620 47780
rect 87780 47420 87800 47780
rect 87460 47400 87800 47420
rect 80400 47300 80800 47320
rect 68900 46200 68960 47220
rect 71900 46300 71960 47280
rect 74400 46400 74460 47280
rect 80220 46500 80280 47240
rect 83120 46600 83180 47280
rect 85620 46700 85680 47280
rect 87240 46800 87300 47280
rect 87240 46740 87900 46800
rect 85620 46640 87900 46700
rect 83120 46540 87900 46600
rect 80220 46440 87900 46500
rect 74400 46340 87900 46400
rect 71900 46240 87900 46300
rect 68900 46140 87900 46200
rect 65200 46040 87900 46100
rect 65200 39820 65260 46040
rect 65740 45940 87900 46000
rect 65740 39820 65800 45940
rect 66440 45840 87900 45900
rect 66440 39820 66500 45840
rect 66980 45740 87900 45800
rect 66980 39820 67040 45740
rect 67680 45640 87900 45700
rect 67680 39820 67740 45640
rect 68220 45540 87900 45600
rect 68220 39820 68280 45540
rect 68920 45440 87900 45500
rect 68920 39820 68980 45440
rect 69460 45340 87900 45400
rect 69460 39820 69520 45340
rect 70160 45240 87900 45300
rect 70160 39820 70220 45240
rect 70700 45140 87900 45200
rect 70700 39820 70760 45140
rect 65200 39800 65280 39820
rect 65200 39660 65210 39800
rect 65270 39660 65280 39800
rect 64880 39540 64980 39650
rect 64880 39340 64980 39460
rect 65200 39404 65280 39660
rect 65740 39790 65820 39820
rect 65740 39660 65750 39790
rect 65810 39660 65820 39790
rect 65400 39540 65600 39640
rect 65200 39290 65223 39404
rect 65257 39290 65280 39404
rect 65400 39340 65600 39460
rect 65740 39404 65820 39660
rect 66440 39790 66520 39820
rect 66440 39660 66450 39790
rect 66510 39660 66520 39790
rect 66020 39540 66220 39640
rect 65200 39260 65280 39290
rect 65740 39290 65763 39404
rect 65797 39290 65820 39404
rect 66020 39360 66220 39460
rect 66440 39404 66520 39660
rect 66980 39790 67060 39820
rect 66980 39660 66990 39790
rect 67050 39660 67060 39790
rect 66640 39540 66840 39640
rect 65740 39260 65820 39290
rect 66440 39290 66463 39404
rect 66497 39290 66520 39404
rect 66640 39360 66840 39460
rect 66980 39404 67060 39660
rect 67680 39790 67760 39820
rect 67680 39670 67690 39790
rect 67750 39670 67760 39790
rect 67260 39540 67460 39640
rect 66440 39260 66520 39290
rect 66980 39290 67003 39404
rect 67037 39290 67060 39404
rect 67260 39360 67460 39460
rect 67680 39404 67760 39670
rect 68220 39800 68300 39820
rect 68220 39680 68230 39800
rect 68290 39680 68300 39800
rect 67880 39540 68080 39640
rect 66980 39260 67060 39290
rect 67680 39290 67703 39404
rect 67737 39290 67760 39404
rect 67880 39360 68080 39460
rect 68220 39404 68300 39680
rect 68920 39790 69000 39820
rect 68920 39670 68930 39790
rect 68990 39670 69000 39790
rect 68500 39540 68700 39640
rect 67680 39260 67760 39290
rect 68220 39290 68243 39404
rect 68277 39290 68300 39404
rect 68500 39360 68700 39460
rect 68920 39404 69000 39670
rect 69460 39790 69540 39820
rect 69460 39670 69470 39790
rect 69530 39670 69540 39790
rect 69120 39540 69320 39640
rect 68220 39260 68300 39290
rect 68920 39290 68943 39404
rect 68977 39290 69000 39404
rect 69120 39360 69320 39460
rect 69460 39404 69540 39670
rect 70160 39790 70240 39820
rect 70160 39670 70170 39790
rect 70230 39670 70240 39790
rect 69740 39540 69940 39640
rect 68920 39260 69000 39290
rect 69460 39290 69483 39404
rect 69517 39290 69540 39404
rect 69740 39360 69940 39460
rect 70160 39404 70240 39670
rect 70700 39790 70780 39820
rect 70700 39670 70710 39790
rect 70770 39670 70780 39790
rect 70360 39540 70560 39640
rect 69460 39260 69540 39290
rect 70160 39290 70183 39404
rect 70217 39290 70240 39404
rect 70360 39360 70560 39460
rect 70700 39404 70780 39670
rect 71000 39540 71100 39640
rect 70160 39260 70240 39290
rect 70700 39290 70723 39404
rect 70757 39290 70780 39404
rect 71000 39360 71100 39460
rect 70700 39260 70780 39290
rect 65140 37030 65340 37040
rect 64880 36860 64980 36970
rect 65140 36950 65160 37030
rect 65320 36950 65340 37030
rect 65690 37030 65880 37050
rect 65140 36900 65340 36950
rect 65200 36850 65280 36900
rect 65400 36870 65600 36970
rect 65690 36950 65700 37030
rect 65860 36950 65880 37030
rect 66380 37030 66570 37050
rect 65690 36920 65880 36950
rect 65200 36710 65210 36850
rect 65270 36710 65280 36850
rect 65200 36650 65280 36710
rect 65740 36850 65820 36920
rect 66020 36870 66220 36970
rect 66380 36950 66390 37030
rect 66560 36950 66570 37030
rect 66930 37030 67120 37050
rect 66380 36930 66570 36950
rect 65740 36720 65750 36850
rect 65810 36720 65820 36850
rect 65740 36650 65820 36720
rect 66440 36850 66520 36930
rect 66640 36870 66840 36970
rect 66930 36950 66940 37030
rect 67100 36950 67120 37030
rect 67610 37030 67820 37060
rect 66930 36930 67120 36950
rect 66440 36720 66450 36850
rect 66510 36720 66520 36850
rect 66440 36650 66520 36720
rect 66980 36850 67060 36930
rect 67260 36870 67460 36970
rect 67610 36950 67630 37030
rect 67800 36950 67820 37030
rect 68160 37030 68350 37050
rect 67610 36930 67820 36950
rect 66980 36720 66990 36850
rect 67050 36720 67060 36850
rect 66980 36650 67060 36720
rect 67680 36840 67760 36930
rect 67880 36870 68080 36970
rect 68160 36950 68180 37030
rect 68340 36950 68350 37030
rect 68860 37030 69040 37050
rect 68160 36930 68350 36950
rect 67680 36720 67690 36840
rect 67750 36720 67760 36840
rect 67680 36650 67760 36720
rect 68220 36830 68300 36930
rect 68500 36870 68700 36970
rect 68860 36950 68880 37030
rect 69020 36950 69040 37030
rect 69400 37030 69600 37050
rect 68860 36930 69040 36950
rect 68220 36710 68230 36830
rect 68290 36710 68300 36830
rect 68220 36650 68300 36710
rect 68920 36840 69000 36930
rect 69120 36870 69320 36970
rect 69400 36950 69420 37030
rect 69580 36950 69600 37030
rect 70100 37030 70300 37050
rect 69400 36930 69600 36950
rect 68920 36720 68930 36840
rect 68990 36720 69000 36840
rect 68920 36650 69000 36720
rect 69460 36840 69540 36930
rect 69740 36870 69940 36970
rect 70100 36950 70120 37030
rect 70280 36950 70300 37030
rect 70640 37030 70840 37050
rect 70100 36930 70300 36950
rect 69460 36720 69470 36840
rect 69530 36720 69540 36840
rect 69460 36650 69540 36720
rect 70160 36840 70240 36930
rect 70360 36870 70560 36970
rect 70640 36950 70660 37030
rect 70820 36950 70840 37030
rect 70640 36930 70840 36950
rect 70160 36720 70170 36840
rect 70230 36720 70240 36840
rect 70160 36650 70240 36720
rect 70700 36840 70780 36930
rect 71000 36870 71100 36970
rect 70700 36720 70710 36840
rect 70770 36720 70780 36840
rect 70700 36650 70780 36720
rect 52080 36580 52400 36600
rect -13400 36180 -13060 36380
rect -13400 35820 -13380 36180
rect -13220 35820 -13060 36180
rect -13400 35800 -13060 35820
rect -600 36180 -260 36380
rect -600 35820 -580 36180
rect -420 35820 -260 36180
rect -600 35800 -260 35820
rect 24800 36180 25240 36380
rect 24800 35820 24820 36180
rect 24980 35820 25240 36180
rect 24800 35800 25240 35820
rect 37600 36180 38040 36380
rect 37600 35820 37620 36180
rect 37780 35820 38040 36180
rect 37600 35800 38040 35820
rect 46720 36180 47000 36380
rect 46720 35820 46820 36180
rect 46980 35820 47000 36180
rect 46720 35800 47000 35820
rect 50080 36180 50400 36380
rect 52080 36220 52220 36580
rect 52380 36220 52400 36580
rect 63240 36580 63600 36600
rect 52080 36200 52400 36220
rect 50080 35820 50220 36180
rect 50380 35820 50400 36180
rect 57920 36180 58200 36380
rect 50080 35800 50400 35820
rect -12200 34060 -12140 35240
rect 600 34160 660 35240
rect 26100 34260 26160 35240
rect 38900 34360 38960 35220
rect 46180 34460 46240 35220
rect 49520 34560 49580 35220
rect 51900 34660 51960 36160
rect 57920 35820 58020 36180
rect 58180 35820 58200 36180
rect 57920 35800 58200 35820
rect 61280 36180 61600 36380
rect 63240 36220 63420 36580
rect 63580 36220 63600 36580
rect 63240 36200 63600 36220
rect 61280 35820 61420 36180
rect 61580 35820 61600 36180
rect 61280 35800 61600 35820
rect 57360 34760 57420 35220
rect 60720 34860 60780 35220
rect 63100 34960 63160 36120
rect 65210 34960 65270 36650
rect 63100 34900 65270 34960
rect 65750 34860 65810 36650
rect 60720 34800 65810 34860
rect 66440 34760 66500 36650
rect 57360 34700 66500 34760
rect 66990 34660 67050 36650
rect 51900 34600 67050 34660
rect 67680 34560 67740 36650
rect 49520 34500 67740 34560
rect 68230 34460 68290 36650
rect 46180 34400 68290 34460
rect 68930 34360 68990 36650
rect 38900 34300 68990 34360
rect 69470 34260 69530 36650
rect 26100 34200 69530 34260
rect 70170 34160 70230 36650
rect 600 34100 70230 34160
rect 70710 34060 70770 36650
rect -12200 34000 70770 34060
<< via1 >>
rect -13380 67420 -13220 67780
rect -580 67420 -420 67780
rect 24820 67420 24980 67780
rect 37620 67420 37780 67780
rect 46820 67420 46980 67780
rect 50220 67420 50380 67780
rect 58020 67420 58180 67780
rect 52220 67020 52380 67380
rect 61420 67420 61580 67780
rect 63420 67020 63580 67380
rect -13800 66480 -13600 66640
rect -13120 66480 -12920 66640
rect -12380 66480 -12180 66640
rect -11540 66380 -11340 66540
rect -10740 66380 -10540 66540
rect -1000 66480 -820 66640
rect -300 66480 -120 66640
rect 440 66480 620 66640
rect 1220 66400 1400 66540
rect 2060 66400 2240 66540
rect 24500 66480 24700 66640
rect 25200 66480 25400 66640
rect 25920 66480 26120 66640
rect 26760 66380 26960 66540
rect 27560 66380 27760 66540
rect 37300 66480 37500 66640
rect 38000 66480 38200 66640
rect 38720 66480 38920 66640
rect 39560 66380 39760 66540
rect 40360 66380 40560 66540
rect 45340 66420 45540 66560
rect 46180 66420 46380 66640
rect 46860 66420 47060 66640
rect 48720 66420 48920 66560
rect 49540 66420 49740 66640
rect 50180 66420 50380 66640
rect 51910 66530 52070 66730
rect 56540 66420 56740 66560
rect 57380 66420 57580 66640
rect 58060 66420 58260 66640
rect 59920 66420 60120 66560
rect 60740 66420 60940 66620
rect 61380 66420 61580 66620
rect 63110 66530 63270 66730
rect 69220 55820 69380 56080
rect 72220 55820 72380 56080
rect 74720 55820 74880 56080
rect 80520 55820 80680 56080
rect 83420 55820 83580 56080
rect 85920 55820 86080 56080
rect 87520 55820 87680 56080
rect 68930 55330 69150 55530
rect 71790 55300 71990 55440
rect 74310 55300 74390 55440
rect 80220 55330 80420 55530
rect 82970 55300 83170 55440
rect 85510 55300 85590 55440
rect 87110 55300 87190 55440
rect 68930 47980 69150 48170
rect 71790 48060 72010 48200
rect 74310 48060 74390 48200
rect 80220 47970 80430 48170
rect 83000 48060 83200 48200
rect 85510 48060 85590 48200
rect 87110 48060 87190 48200
rect 69220 47320 69380 47680
rect 72220 47420 72380 47780
rect 74720 47420 74880 47780
rect 80620 47320 80780 47680
rect 83420 47420 83580 47780
rect 86020 47420 86180 47780
rect 87620 47420 87780 47780
rect 65430 38310 65590 38490
rect 66670 38310 66830 38490
rect 67910 38310 68070 38490
rect 69150 38310 69310 38490
rect 70390 38310 70550 38490
rect 65430 37310 65590 37490
rect 66670 37310 66830 37490
rect 67910 37310 68070 37490
rect 69150 37310 69310 37490
rect 70390 37310 70550 37490
rect -13800 36960 -13560 37120
rect -13100 36960 -12860 37120
rect -12420 36960 -12180 37120
rect -11560 37060 -11320 37220
rect -10780 37060 -10540 37220
rect -1000 36960 -760 37120
rect -360 36960 -120 37120
rect 380 36960 620 37120
rect 1240 37060 1480 37220
rect 2020 37060 2260 37220
rect 24500 36960 24800 37120
rect 25140 36960 25440 37120
rect 25820 36960 26120 37120
rect 26660 37060 26960 37220
rect 27460 37060 27760 37220
rect 37300 36960 37600 37120
rect 37960 36960 38260 37120
rect 38620 36960 38920 37120
rect 39440 37060 39740 37220
rect 40260 37060 40560 37220
rect 45340 37040 45580 37180
rect 46180 36960 46420 37180
rect 46820 36960 47060 37180
rect 48720 37040 49000 37180
rect 49540 36960 49820 37180
rect 50100 36960 50380 37180
rect 51910 36870 52070 37070
rect 56540 37040 56780 37180
rect 57380 36960 57580 37180
rect 58060 36960 58260 37180
rect 59920 37040 60100 37180
rect 60740 36960 60920 37180
rect 61400 36960 61580 37180
rect 63120 36880 63260 37060
rect -13380 35820 -13220 36180
rect -580 35820 -420 36180
rect 24820 35820 24980 36180
rect 37620 35820 37780 36180
rect 46820 35820 46980 36180
rect 52220 36220 52380 36580
rect 50220 35820 50380 36180
rect 58020 35820 58180 36180
rect 63420 36220 63580 36580
rect 61420 35820 61580 36180
<< metal2 >>
rect -13400 67780 -13200 67800
rect -13400 67420 -13380 67780
rect -13220 67420 -13200 67780
rect -13400 67400 -13200 67420
rect -600 67780 -400 67800
rect -600 67420 -580 67780
rect -420 67420 -400 67780
rect -600 67400 -400 67420
rect 24800 67780 25000 67800
rect 24800 67420 24820 67780
rect 24980 67420 25000 67780
rect 24800 67400 25000 67420
rect 37600 67780 37800 67800
rect 37600 67420 37620 67780
rect 37780 67420 37800 67780
rect 37600 67400 37800 67420
rect 46800 67780 47000 67800
rect 46800 67420 46820 67780
rect 46980 67420 47000 67780
rect 46800 67400 47000 67420
rect 50200 67780 50400 67800
rect 50200 67420 50220 67780
rect 50380 67420 50400 67780
rect 50200 67400 50400 67420
rect 58000 67780 58200 67800
rect 58000 67420 58020 67780
rect 58180 67420 58200 67780
rect 58000 67400 58200 67420
rect 61400 67780 61600 67800
rect 61400 67420 61420 67780
rect 61580 67420 61600 67780
rect 61400 67400 61600 67420
rect 52200 67380 52400 67400
rect 52200 67020 52220 67380
rect 52380 67020 52400 67380
rect 52200 67000 52400 67020
rect 63400 67380 63600 67400
rect 63400 67020 63420 67380
rect 63580 67020 63600 67380
rect 63400 67000 63600 67020
rect 51900 66730 52080 66740
rect -13820 66640 -13580 66660
rect -13820 66480 -13800 66640
rect -13600 66480 -13580 66640
rect -13820 66180 -13580 66480
rect -13820 65920 -13800 66180
rect -13600 65920 -13580 66180
rect -13820 65900 -13580 65920
rect -13140 66640 -12900 66660
rect -13140 66480 -13120 66640
rect -12920 66480 -12900 66640
rect -13140 66180 -12900 66480
rect -13140 65920 -13120 66180
rect -12920 65920 -12900 66180
rect -13140 65900 -12900 65920
rect -12400 66640 -12160 66660
rect -12400 66480 -12380 66640
rect -12180 66480 -12160 66640
rect -1020 66640 -800 66660
rect -12400 66180 -12160 66480
rect -12400 65920 -12380 66180
rect -12180 65920 -12160 66180
rect -12400 65900 -12160 65920
rect -11560 66540 -11320 66560
rect -11560 66380 -11540 66540
rect -11340 66380 -11320 66540
rect -11560 66180 -11320 66380
rect -11560 65920 -11540 66180
rect -11340 65920 -11320 66180
rect -11560 65900 -11320 65920
rect -10760 66540 -10520 66560
rect -10760 66380 -10740 66540
rect -10540 66380 -10520 66540
rect -10760 66180 -10520 66380
rect -10760 65920 -10740 66180
rect -10540 65920 -10520 66180
rect -10760 65900 -10520 65920
rect -1020 66480 -1000 66640
rect -820 66480 -800 66640
rect -1020 66180 -800 66480
rect -1020 65920 -1000 66180
rect -820 65920 -800 66180
rect -1020 65900 -800 65920
rect -320 66640 -100 66660
rect -320 66480 -300 66640
rect -120 66480 -100 66640
rect -320 66180 -100 66480
rect -320 65920 -300 66180
rect -120 65920 -100 66180
rect -320 65900 -100 65920
rect 420 66640 640 66660
rect 420 66480 440 66640
rect 620 66480 640 66640
rect 24480 66640 24720 66660
rect 420 66180 640 66480
rect 420 65920 440 66180
rect 620 65920 640 66180
rect 420 65900 640 65920
rect 1200 66540 1420 66560
rect 1200 66400 1220 66540
rect 1400 66400 1420 66540
rect 1200 66180 1420 66400
rect 1200 65920 1220 66180
rect 1400 65920 1420 66180
rect 1200 65900 1420 65920
rect 2040 66540 2260 66560
rect 2040 66400 2060 66540
rect 2240 66400 2260 66540
rect 2040 66180 2260 66400
rect 2040 65920 2060 66180
rect 2240 65920 2260 66180
rect 2040 65900 2260 65920
rect 24480 66480 24500 66640
rect 24700 66480 24720 66640
rect 24480 66180 24720 66480
rect 24480 65920 24500 66180
rect 24700 65920 24720 66180
rect 24480 65900 24720 65920
rect 25180 66640 25420 66660
rect 25180 66480 25200 66640
rect 25400 66480 25420 66640
rect 25180 66180 25420 66480
rect 25180 65920 25200 66180
rect 25400 65920 25420 66180
rect 25180 65900 25420 65920
rect 25900 66640 26140 66660
rect 25900 66480 25920 66640
rect 26120 66480 26140 66640
rect 37280 66640 37520 66660
rect 25900 66180 26140 66480
rect 25900 65920 25920 66180
rect 26120 65920 26140 66180
rect 25900 65900 26140 65920
rect 26740 66540 26980 66560
rect 26740 66380 26760 66540
rect 26960 66380 26980 66540
rect 26740 66180 26980 66380
rect 26740 65920 26760 66180
rect 26960 65920 26980 66180
rect 26740 65900 26980 65920
rect 27540 66540 27780 66560
rect 27540 66380 27560 66540
rect 27760 66380 27780 66540
rect 27540 66180 27780 66380
rect 27540 65920 27560 66180
rect 27760 65920 27780 66180
rect 27540 65900 27780 65920
rect 37280 66480 37300 66640
rect 37500 66480 37520 66640
rect 37280 66180 37520 66480
rect 37280 65920 37300 66180
rect 37500 65920 37520 66180
rect 37280 65900 37520 65920
rect 37980 66640 38220 66660
rect 37980 66480 38000 66640
rect 38200 66480 38220 66640
rect 37980 66180 38220 66480
rect 37980 65920 38000 66180
rect 38200 65920 38220 66180
rect 37980 65900 38220 65920
rect 38700 66640 38940 66660
rect 38700 66480 38720 66640
rect 38920 66480 38940 66640
rect 46160 66640 46400 66660
rect 45320 66560 45560 66580
rect 38700 66180 38940 66480
rect 38700 65920 38720 66180
rect 38920 65920 38940 66180
rect 38700 65900 38940 65920
rect 39540 66540 39780 66560
rect 39540 66380 39560 66540
rect 39760 66380 39780 66540
rect 39540 66180 39780 66380
rect 39540 65920 39560 66180
rect 39760 65920 39780 66180
rect 39540 65900 39780 65920
rect 40340 66540 40580 66560
rect 40340 66380 40360 66540
rect 40560 66380 40580 66540
rect 40340 66180 40580 66380
rect 40340 65920 40360 66180
rect 40560 65920 40580 66180
rect 40340 65900 40580 65920
rect 45320 66420 45340 66560
rect 45540 66420 45560 66560
rect 45320 66180 45560 66420
rect 45320 65920 45340 66180
rect 45540 65920 45560 66180
rect 45320 65900 45560 65920
rect 46160 66420 46180 66640
rect 46380 66420 46400 66640
rect 46160 66180 46400 66420
rect 46160 65920 46180 66180
rect 46380 65920 46400 66180
rect 46160 65900 46400 65920
rect 46840 66640 47080 66660
rect 46840 66420 46860 66640
rect 47060 66420 47080 66640
rect 49520 66640 49760 66660
rect 46840 66180 47080 66420
rect 46840 65920 46860 66180
rect 47060 65920 47080 66180
rect 46840 65900 47080 65920
rect 48700 66560 48940 66580
rect 48700 66420 48720 66560
rect 48920 66420 48940 66560
rect 48700 66180 48940 66420
rect 48700 65920 48720 66180
rect 48920 65920 48940 66180
rect 48700 65900 48940 65920
rect 49520 66420 49540 66640
rect 49740 66420 49760 66640
rect 49520 66180 49760 66420
rect 49520 65920 49540 66180
rect 49740 65920 49760 66180
rect 49520 65900 49760 65920
rect 50160 66640 50400 66660
rect 50160 66420 50180 66640
rect 50380 66420 50400 66640
rect 50160 66180 50400 66420
rect 50160 65920 50180 66180
rect 50380 65920 50400 66180
rect 50160 65900 50400 65920
rect 51900 66530 51910 66730
rect 52070 66530 52080 66730
rect 63100 66730 63280 66740
rect 57360 66640 57600 66660
rect 51900 66190 52080 66530
rect 51900 65920 51910 66190
rect 52070 65920 52080 66190
rect 51900 65910 52080 65920
rect 56520 66560 56760 66580
rect 56520 66420 56540 66560
rect 56740 66420 56760 66560
rect 56520 66180 56760 66420
rect 56520 65920 56540 66180
rect 56740 65920 56760 66180
rect 56520 65900 56760 65920
rect 57360 66420 57380 66640
rect 57580 66420 57600 66640
rect 57360 66180 57600 66420
rect 57360 65920 57380 66180
rect 57580 65920 57600 66180
rect 57360 65900 57600 65920
rect 58040 66640 58280 66660
rect 58040 66420 58060 66640
rect 58260 66420 58280 66640
rect 60720 66620 60960 66640
rect 58040 66180 58280 66420
rect 58040 65920 58060 66180
rect 58260 65920 58280 66180
rect 58040 65900 58280 65920
rect 59900 66560 60140 66580
rect 59900 66420 59920 66560
rect 60120 66420 60140 66560
rect 59900 66180 60140 66420
rect 59900 65920 59920 66180
rect 60120 65920 60140 66180
rect 59900 65900 60140 65920
rect 60720 66420 60740 66620
rect 60940 66420 60960 66620
rect 60720 66180 60960 66420
rect 60720 65920 60740 66180
rect 60940 65920 60960 66180
rect 60720 65900 60960 65920
rect 61360 66620 61600 66640
rect 61360 66420 61380 66620
rect 61580 66420 61600 66620
rect 61360 66180 61600 66420
rect 61360 65920 61380 66180
rect 61580 65920 61600 66180
rect 61360 65900 61600 65920
rect 63100 66530 63110 66730
rect 63270 66530 63280 66730
rect 63100 66190 63280 66530
rect 63100 65920 63110 66190
rect 63270 65920 63280 66190
rect 63100 65910 63280 65920
rect 69200 56080 69400 56100
rect 69200 55820 69220 56080
rect 69380 55820 69400 56080
rect 69200 55800 69400 55820
rect 72200 56080 72400 56100
rect 72200 55820 72220 56080
rect 72380 55820 72400 56080
rect 72200 55800 72400 55820
rect 74700 56080 74900 56100
rect 74700 55820 74720 56080
rect 74880 55820 74900 56080
rect 74700 55800 74900 55820
rect 80500 56080 80700 56100
rect 80500 55820 80520 56080
rect 80680 55820 80700 56080
rect 80500 55800 80700 55820
rect 83400 56080 83600 56100
rect 83400 55820 83420 56080
rect 83580 55820 83600 56080
rect 83400 55800 83600 55820
rect 85900 56080 86100 56100
rect 85900 55820 85920 56080
rect 86080 55820 86100 56080
rect 85900 55800 86100 55820
rect 87500 56080 87700 56100
rect 87500 55820 87520 56080
rect 87680 55820 87700 56080
rect 87500 55800 87700 55820
rect 68920 55530 69160 55540
rect 68920 55330 68930 55530
rect 69150 55330 69160 55530
rect 80210 55530 80430 55540
rect 68920 54990 69160 55330
rect 68920 54710 68930 54990
rect 69150 54710 69160 54990
rect 68920 54700 69160 54710
rect 71780 55440 72000 55450
rect 71780 55300 71790 55440
rect 71990 55300 72000 55440
rect 71780 54990 72000 55300
rect 71780 54710 71790 54990
rect 71990 54710 72000 54990
rect 74300 55440 74400 55450
rect 74300 55300 74310 55440
rect 74390 55300 74400 55440
rect 74300 54990 74400 55300
rect 74300 54770 74310 54990
rect 74390 54770 74400 54990
rect 74300 54760 74400 54770
rect 80210 55330 80220 55530
rect 80420 55330 80430 55530
rect 80210 54990 80430 55330
rect 71780 54700 72000 54710
rect 80210 54710 80220 54990
rect 80420 54710 80430 54990
rect 80210 54700 80430 54710
rect 82960 55440 83180 55450
rect 82960 55300 82970 55440
rect 83170 55300 83180 55440
rect 82960 54990 83180 55300
rect 82960 54710 82970 54990
rect 83170 54710 83180 54990
rect 85500 55440 85600 55450
rect 85500 55300 85510 55440
rect 85590 55300 85600 55440
rect 85500 54990 85600 55300
rect 85500 54770 85510 54990
rect 85590 54770 85600 54990
rect 85500 54760 85600 54770
rect 87100 55440 87200 55450
rect 87100 55300 87110 55440
rect 87190 55300 87200 55440
rect 87100 54990 87200 55300
rect 87100 54770 87110 54990
rect 87190 54770 87200 54990
rect 87100 54760 87200 54770
rect 82960 54700 83180 54710
rect 68920 48890 69160 48900
rect 68920 48610 68930 48890
rect 69150 48610 69160 48890
rect 68920 48170 69160 48610
rect 68920 47980 68930 48170
rect 69150 47980 69160 48170
rect 71780 48890 72020 48900
rect 71780 48610 71790 48890
rect 72010 48610 72020 48890
rect 80210 48890 80440 48900
rect 71780 48200 72020 48610
rect 71780 48060 71790 48200
rect 72010 48060 72020 48200
rect 71780 48050 72020 48060
rect 74300 48830 74400 48840
rect 74300 48610 74310 48830
rect 74390 48610 74400 48830
rect 74300 48200 74400 48610
rect 74300 48060 74310 48200
rect 74390 48060 74400 48200
rect 74300 48050 74400 48060
rect 80210 48610 80220 48890
rect 80430 48610 80440 48890
rect 80210 48170 80440 48610
rect 68920 47970 69160 47980
rect 80210 47970 80220 48170
rect 80430 47970 80440 48170
rect 82990 48890 83210 48900
rect 82990 48610 83000 48890
rect 83200 48610 83210 48890
rect 82990 48200 83210 48610
rect 82990 48060 83000 48200
rect 83200 48060 83210 48200
rect 82990 48050 83210 48060
rect 85500 48870 85600 48880
rect 85500 48610 85510 48870
rect 85590 48610 85600 48870
rect 85500 48200 85600 48610
rect 85500 48060 85510 48200
rect 85590 48060 85600 48200
rect 85500 48050 85600 48060
rect 87100 48870 87200 48880
rect 87100 48610 87110 48870
rect 87190 48610 87200 48870
rect 87100 48200 87200 48610
rect 87100 48060 87110 48200
rect 87190 48060 87200 48200
rect 87100 48050 87200 48060
rect 80210 47960 80440 47970
rect 72200 47780 72400 47800
rect 69200 47680 69400 47700
rect 69200 47320 69220 47680
rect 69380 47320 69400 47680
rect 72200 47420 72220 47780
rect 72380 47420 72400 47780
rect 72200 47400 72400 47420
rect 74700 47780 74900 47800
rect 74700 47420 74720 47780
rect 74880 47420 74900 47780
rect 83400 47780 83600 47800
rect 74700 47400 74900 47420
rect 80600 47680 80800 47700
rect 69200 47200 69400 47320
rect 80600 47320 80620 47680
rect 80780 47320 80800 47680
rect 83400 47420 83420 47780
rect 83580 47420 83600 47780
rect 83400 47400 83600 47420
rect 86000 47780 86200 47800
rect 86000 47420 86020 47780
rect 86180 47420 86200 47780
rect 86000 47400 86200 47420
rect 87600 47780 87800 47800
rect 87600 47420 87620 47780
rect 87780 47420 87800 47780
rect 87600 47400 87800 47420
rect 80600 47200 80800 47320
rect 65420 38490 65600 38500
rect 65420 38310 65430 38490
rect 65590 38310 65600 38490
rect 65420 38300 65600 38310
rect 66660 38490 66840 38500
rect 66660 38310 66670 38490
rect 66830 38310 66840 38490
rect 66660 38300 66840 38310
rect 67900 38490 68080 38500
rect 67900 38310 67910 38490
rect 68070 38310 68080 38490
rect 67900 38300 68080 38310
rect 69140 38490 69320 38500
rect 69140 38310 69150 38490
rect 69310 38310 69320 38490
rect 69140 38300 69320 38310
rect 70380 38490 70560 38500
rect 70380 38310 70390 38490
rect 70550 38310 70560 38490
rect 70380 38300 70560 38310
rect -13820 37680 -13540 37700
rect -13820 37420 -13800 37680
rect -13560 37420 -13540 37680
rect -13820 37120 -13540 37420
rect -13820 36960 -13800 37120
rect -13560 36960 -13540 37120
rect -13820 36940 -13540 36960
rect -13120 37680 -12840 37700
rect -13120 37420 -13100 37680
rect -12860 37420 -12840 37680
rect -13120 37120 -12840 37420
rect -13120 36960 -13100 37120
rect -12860 36960 -12840 37120
rect -13120 36940 -12840 36960
rect -12440 37680 -12160 37700
rect -12440 37420 -12420 37680
rect -12180 37420 -12160 37680
rect -12440 37120 -12160 37420
rect -12440 36960 -12420 37120
rect -12180 36960 -12160 37120
rect -11580 37680 -11300 37700
rect -11580 37420 -11560 37680
rect -11320 37420 -11300 37680
rect -11580 37220 -11300 37420
rect -11580 37060 -11560 37220
rect -11320 37060 -11300 37220
rect -11580 37040 -11300 37060
rect -10800 37680 -10520 37700
rect -10800 37420 -10780 37680
rect -10540 37420 -10520 37680
rect -10800 37220 -10520 37420
rect -10800 37060 -10780 37220
rect -10540 37060 -10520 37220
rect -10800 37040 -10520 37060
rect -1020 37680 -740 37700
rect -1020 37420 -1000 37680
rect -760 37420 -740 37680
rect -1020 37120 -740 37420
rect -12440 36940 -12160 36960
rect -1020 36960 -1000 37120
rect -760 36960 -740 37120
rect -1020 36940 -740 36960
rect -380 37680 -100 37700
rect -380 37420 -360 37680
rect -120 37420 -100 37680
rect -380 37120 -100 37420
rect -380 36960 -360 37120
rect -120 36960 -100 37120
rect -380 36940 -100 36960
rect 360 37680 640 37700
rect 360 37420 380 37680
rect 620 37420 640 37680
rect 360 37120 640 37420
rect 360 36960 380 37120
rect 620 36960 640 37120
rect 1220 37680 1500 37700
rect 1220 37420 1240 37680
rect 1480 37420 1500 37680
rect 1220 37220 1500 37420
rect 1220 37060 1240 37220
rect 1480 37060 1500 37220
rect 1220 37040 1500 37060
rect 2000 37680 2280 37700
rect 2000 37420 2020 37680
rect 2260 37420 2280 37680
rect 2000 37220 2280 37420
rect 2000 37060 2020 37220
rect 2260 37060 2280 37220
rect 2000 37040 2280 37060
rect 24480 37680 24820 37700
rect 24480 37420 24500 37680
rect 24800 37420 24820 37680
rect 24480 37120 24820 37420
rect 360 36940 640 36960
rect 24480 36960 24500 37120
rect 24800 36960 24820 37120
rect 24480 36940 24820 36960
rect 25120 37680 25460 37700
rect 25120 37420 25140 37680
rect 25440 37420 25460 37680
rect 25120 37120 25460 37420
rect 25120 36960 25140 37120
rect 25440 36960 25460 37120
rect 25120 36940 25460 36960
rect 25800 37680 26140 37700
rect 25800 37420 25820 37680
rect 26120 37420 26140 37680
rect 25800 37120 26140 37420
rect 25800 36960 25820 37120
rect 26120 36960 26140 37120
rect 26640 37680 26980 37700
rect 26640 37420 26660 37680
rect 26960 37420 26980 37680
rect 26640 37220 26980 37420
rect 26640 37060 26660 37220
rect 26960 37060 26980 37220
rect 26640 37040 26980 37060
rect 27440 37680 27780 37700
rect 27440 37420 27460 37680
rect 27760 37420 27780 37680
rect 27440 37220 27780 37420
rect 27440 37060 27460 37220
rect 27760 37060 27780 37220
rect 27440 37040 27780 37060
rect 37280 37680 37620 37700
rect 37280 37420 37300 37680
rect 37600 37420 37620 37680
rect 37280 37120 37620 37420
rect 25800 36940 26140 36960
rect 37280 36960 37300 37120
rect 37600 36960 37620 37120
rect 37280 36940 37620 36960
rect 37940 37680 38280 37700
rect 37940 37420 37960 37680
rect 38260 37420 38280 37680
rect 37940 37120 38280 37420
rect 37940 36960 37960 37120
rect 38260 36960 38280 37120
rect 37940 36940 38280 36960
rect 38600 37680 38940 37700
rect 38600 37420 38620 37680
rect 38920 37420 38940 37680
rect 38600 37120 38940 37420
rect 38600 36960 38620 37120
rect 38920 36960 38940 37120
rect 39420 37680 39760 37700
rect 39420 37420 39440 37680
rect 39740 37420 39760 37680
rect 39420 37220 39760 37420
rect 39420 37060 39440 37220
rect 39740 37060 39760 37220
rect 39420 37040 39760 37060
rect 40240 37680 40580 37700
rect 40240 37420 40260 37680
rect 40560 37420 40580 37680
rect 40240 37220 40580 37420
rect 40240 37060 40260 37220
rect 40560 37060 40580 37220
rect 40240 37040 40580 37060
rect 45320 37680 45600 37700
rect 45320 37420 45340 37680
rect 45580 37420 45600 37680
rect 45320 37180 45600 37420
rect 45320 37040 45340 37180
rect 45580 37040 45600 37180
rect 45320 37020 45600 37040
rect 46160 37680 46440 37700
rect 46160 37420 46180 37680
rect 46420 37420 46440 37680
rect 46160 37180 46440 37420
rect 38600 36940 38940 36960
rect 46160 36960 46180 37180
rect 46420 36960 46440 37180
rect 46160 36940 46440 36960
rect 46800 37680 47080 37700
rect 46800 37420 46820 37680
rect 47060 37420 47080 37680
rect 46800 37180 47080 37420
rect 46800 36960 46820 37180
rect 47060 36960 47080 37180
rect 48700 37680 49020 37700
rect 48700 37420 48720 37680
rect 49000 37420 49020 37680
rect 48700 37180 49020 37420
rect 48700 37040 48720 37180
rect 49000 37040 49020 37180
rect 48700 37020 49020 37040
rect 49520 37680 49840 37700
rect 49520 37420 49540 37680
rect 49820 37420 49840 37680
rect 49520 37180 49840 37420
rect 46800 36940 47080 36960
rect 49520 36960 49540 37180
rect 49820 36960 49840 37180
rect 49520 36940 49840 36960
rect 50080 37680 50400 37700
rect 50080 37420 50100 37680
rect 50380 37420 50400 37680
rect 50080 37180 50400 37420
rect 50080 36960 50100 37180
rect 50380 36960 50400 37180
rect 50080 36940 50400 36960
rect 51900 37680 52080 37700
rect 51900 37420 51920 37680
rect 52060 37420 52080 37680
rect 51900 37070 52080 37420
rect 51900 36870 51910 37070
rect 52070 36870 52080 37070
rect 56520 37680 56800 37700
rect 56520 37420 56540 37680
rect 56780 37420 56800 37680
rect 56520 37180 56800 37420
rect 56520 37040 56540 37180
rect 56780 37040 56800 37180
rect 56520 37020 56800 37040
rect 57360 37680 57600 37700
rect 57360 37420 57380 37680
rect 57580 37420 57600 37680
rect 57360 37180 57600 37420
rect 57360 36960 57380 37180
rect 57580 36960 57600 37180
rect 57360 36940 57600 36960
rect 58040 37680 58280 37700
rect 58040 37420 58060 37680
rect 58260 37420 58280 37680
rect 58040 37180 58280 37420
rect 58040 36960 58060 37180
rect 58260 36960 58280 37180
rect 59900 37680 60120 37700
rect 59900 37420 59920 37680
rect 60100 37420 60120 37680
rect 59900 37180 60120 37420
rect 59900 37040 59920 37180
rect 60100 37040 60120 37180
rect 59900 37020 60120 37040
rect 60720 37680 60940 37700
rect 60720 37420 60740 37680
rect 60920 37420 60940 37680
rect 60720 37180 60940 37420
rect 58040 36940 58280 36960
rect 60720 36960 60740 37180
rect 60920 36960 60940 37180
rect 60720 36940 60940 36960
rect 61380 37680 61600 37700
rect 61380 37420 61400 37680
rect 61580 37420 61600 37680
rect 61380 37180 61600 37420
rect 61380 36960 61400 37180
rect 61580 36960 61600 37180
rect 61380 36940 61600 36960
rect 63100 37640 63280 37660
rect 63100 37420 63120 37640
rect 63260 37420 63280 37640
rect 63100 37060 63280 37420
rect 65420 37490 65600 37500
rect 65420 37310 65430 37490
rect 65590 37310 65600 37490
rect 65420 37300 65600 37310
rect 66660 37490 66840 37500
rect 66660 37310 66670 37490
rect 66830 37310 66840 37490
rect 66660 37300 66840 37310
rect 67900 37490 68080 37500
rect 67900 37310 67910 37490
rect 68070 37310 68080 37490
rect 67900 37300 68080 37310
rect 69140 37490 69320 37500
rect 69140 37310 69150 37490
rect 69310 37310 69320 37490
rect 69140 37300 69320 37310
rect 70380 37490 70560 37500
rect 70380 37310 70390 37490
rect 70550 37310 70560 37490
rect 70380 37300 70560 37310
rect 51900 36860 52080 36870
rect 63100 36880 63120 37060
rect 63260 36880 63280 37060
rect 63100 36860 63280 36880
rect 52200 36580 52400 36600
rect 52200 36220 52220 36580
rect 52380 36220 52400 36580
rect 52200 36200 52400 36220
rect 63400 36580 63600 36600
rect 63400 36220 63420 36580
rect 63580 36220 63600 36580
rect 63400 36200 63600 36220
rect -13400 36180 -13200 36200
rect -13400 35820 -13380 36180
rect -13220 35820 -13200 36180
rect -13400 35800 -13200 35820
rect -600 36180 -400 36200
rect -600 35820 -580 36180
rect -420 35820 -400 36180
rect -600 35800 -400 35820
rect 24800 36180 25000 36200
rect 24800 35820 24820 36180
rect 24980 35820 25000 36180
rect 24800 35800 25000 35820
rect 37600 36180 37800 36200
rect 37600 35820 37620 36180
rect 37780 35820 37800 36180
rect 37600 35800 37800 35820
rect 46800 36180 47000 36200
rect 46800 35820 46820 36180
rect 46980 35820 47000 36180
rect 46800 35800 47000 35820
rect 50200 36180 50400 36200
rect 50200 35820 50220 36180
rect 50380 35820 50400 36180
rect 50200 35800 50400 35820
rect 58000 36180 58200 36200
rect 58000 35820 58020 36180
rect 58180 35820 58200 36180
rect 58000 35800 58200 35820
rect 61400 36180 61600 36200
rect 61400 35820 61420 36180
rect 61580 35820 61600 36180
rect 61400 35800 61600 35820
<< via2 >>
rect -13380 67420 -13220 67780
rect -580 67420 -420 67780
rect 24820 67420 24980 67780
rect 37620 67420 37780 67780
rect 46820 67420 46980 67780
rect 50220 67420 50380 67780
rect 58020 67420 58180 67780
rect 61420 67420 61580 67780
rect 52220 67020 52380 67380
rect 63420 67020 63580 67380
rect -13800 65920 -13600 66180
rect -13120 65920 -12920 66180
rect -12380 65920 -12180 66180
rect -11540 65920 -11340 66180
rect -10740 65920 -10540 66180
rect -1000 65920 -820 66180
rect -300 65920 -120 66180
rect 440 65920 620 66180
rect 1220 65920 1400 66180
rect 2060 65920 2240 66180
rect 24500 65920 24700 66180
rect 25200 65920 25400 66180
rect 25920 65920 26120 66180
rect 26760 65920 26960 66180
rect 27560 65920 27760 66180
rect 37300 65920 37500 66180
rect 38000 65920 38200 66180
rect 38720 65920 38920 66180
rect 39560 65920 39760 66180
rect 40360 65920 40560 66180
rect 45340 65920 45540 66180
rect 46180 65920 46380 66180
rect 46860 65920 47060 66180
rect 48720 65920 48920 66180
rect 49540 65920 49740 66180
rect 50180 65920 50380 66180
rect 51910 65920 52070 66190
rect 56540 65920 56740 66180
rect 57380 65920 57580 66180
rect 58060 65920 58260 66180
rect 59920 65920 60120 66180
rect 60740 65920 60940 66180
rect 61380 65920 61580 66180
rect 63110 65920 63270 66190
rect 69220 55820 69380 56080
rect 72220 55820 72380 56080
rect 74720 55820 74880 56080
rect 80520 55820 80680 56080
rect 83420 55820 83580 56080
rect 85920 55820 86080 56080
rect 87520 55820 87680 56080
rect 68930 54710 69150 54990
rect 71790 54710 71990 54990
rect 74310 54770 74390 54990
rect 80220 54710 80420 54990
rect 82970 54710 83170 54990
rect 85510 54770 85590 54990
rect 87110 54770 87190 54990
rect 68930 48610 69150 48890
rect 71790 48610 72010 48890
rect 74310 48610 74390 48830
rect 80220 48610 80430 48890
rect 83000 48610 83200 48890
rect 85510 48610 85590 48870
rect 87110 48610 87190 48870
rect 69220 47320 69380 47680
rect 72220 47420 72380 47780
rect 74720 47420 74880 47780
rect 80620 47320 80780 47680
rect 83420 47420 83580 47780
rect 86020 47420 86180 47780
rect 87620 47420 87780 47780
rect 65430 38310 65590 38490
rect 66670 38310 66830 38490
rect 67910 38310 68070 38490
rect 69150 38310 69310 38490
rect 70390 38310 70550 38490
rect -13800 37420 -13560 37680
rect -13100 37420 -12860 37680
rect -12420 37420 -12180 37680
rect -11560 37420 -11320 37680
rect -10780 37420 -10540 37680
rect -1000 37420 -760 37680
rect -360 37420 -120 37680
rect 380 37420 620 37680
rect 1240 37420 1480 37680
rect 2020 37420 2260 37680
rect 24500 37420 24800 37680
rect 25140 37420 25440 37680
rect 25820 37420 26120 37680
rect 26660 37420 26960 37680
rect 27460 37420 27760 37680
rect 37300 37420 37600 37680
rect 37960 37420 38260 37680
rect 38620 37420 38920 37680
rect 39440 37420 39740 37680
rect 40260 37420 40560 37680
rect 45340 37420 45580 37680
rect 46180 37420 46420 37680
rect 46820 37420 47060 37680
rect 48720 37420 49000 37680
rect 49540 37420 49820 37680
rect 50100 37420 50380 37680
rect 51920 37420 52060 37680
rect 56540 37420 56780 37680
rect 57380 37420 57580 37680
rect 58060 37420 58260 37680
rect 59920 37420 60100 37680
rect 60740 37420 60920 37680
rect 61400 37420 61580 37680
rect 63120 37420 63260 37640
rect 65430 37310 65590 37490
rect 66670 37310 66830 37490
rect 67910 37310 68070 37490
rect 69150 37310 69310 37490
rect 70390 37310 70550 37490
rect 52220 36220 52380 36580
rect 63420 36220 63580 36580
rect -13380 35820 -13220 36180
rect -580 35820 -420 36180
rect 24820 35820 24980 36180
rect 37620 35820 37780 36180
rect 46820 35820 46980 36180
rect 50220 35820 50380 36180
rect 58020 35820 58180 36180
rect 61420 35820 61580 36180
<< metal3 >>
rect -13400 69900 71700 70300
rect -13400 67780 -13200 69900
rect -13400 67420 -13380 67780
rect -13220 67420 -13200 67780
rect -13400 67400 -13200 67420
rect -600 67780 -400 69900
rect -600 67420 -580 67780
rect -420 67420 -400 67780
rect -600 67400 -400 67420
rect 24800 67780 25000 69900
rect 24800 67420 24820 67780
rect 24980 67420 25000 67780
rect 24800 67400 25000 67420
rect 37600 67780 37800 69900
rect 37600 67420 37620 67780
rect 37780 67420 37800 67780
rect 37600 67400 37800 67420
rect 46800 67780 47000 69900
rect 46800 67420 46820 67780
rect 46980 67420 47000 67780
rect 46800 67400 47000 67420
rect 50200 67780 50400 69900
rect 50200 67420 50220 67780
rect 50380 67420 50400 67780
rect 50200 67400 50400 67420
rect 52200 67380 52400 69900
rect 58000 67780 58200 69900
rect 58000 67420 58020 67780
rect 58180 67420 58200 67780
rect 58000 67400 58200 67420
rect 61400 67780 61600 69900
rect 61400 67420 61420 67780
rect 61580 67420 61600 67780
rect 61400 67400 61600 67420
rect 52200 67020 52220 67380
rect 52380 67020 52400 67380
rect 52200 67000 52400 67020
rect 63400 67380 63600 69900
rect 63400 67020 63420 67380
rect 63580 67020 63600 67380
rect 63400 67000 63600 67020
rect 71300 66200 71700 69900
rect -13820 66180 -13580 66200
rect -13820 65920 -13800 66180
rect -13600 65920 -13580 66180
rect -13820 65900 -13580 65920
rect -13140 66180 -12900 66200
rect -13140 65920 -13120 66180
rect -12920 65920 -12900 66180
rect -13140 65900 -12900 65920
rect -12400 66180 -12160 66200
rect -12400 65920 -12380 66180
rect -12180 65920 -12160 66180
rect -12400 65900 -12160 65920
rect -11560 66180 -11320 66200
rect -11560 65920 -11540 66180
rect -11340 65920 -11320 66180
rect -11560 65900 -11320 65920
rect -10760 66180 -10520 66200
rect -10760 65920 -10740 66180
rect -10540 65920 -10520 66180
rect -10760 65900 -10520 65920
rect -1020 66180 -800 66200
rect -1020 65920 -1000 66180
rect -820 65920 -800 66180
rect -1020 65900 -800 65920
rect -320 66180 -100 66200
rect -320 65920 -300 66180
rect -120 65920 -100 66180
rect -320 65900 -100 65920
rect 420 66180 640 66200
rect 420 65920 440 66180
rect 620 65920 640 66180
rect 420 65900 640 65920
rect 1200 66180 1420 66200
rect 1200 65920 1220 66180
rect 1400 65920 1420 66180
rect 1200 65900 1420 65920
rect 2040 66180 2260 66200
rect 2040 65920 2060 66180
rect 2240 65920 2260 66180
rect 2040 65900 2260 65920
rect 24480 66180 24720 66200
rect 24480 65920 24500 66180
rect 24700 65920 24720 66180
rect 24480 65900 24720 65920
rect 25180 66180 25420 66200
rect 25180 65920 25200 66180
rect 25400 65920 25420 66180
rect 25180 65900 25420 65920
rect 25900 66180 26140 66200
rect 25900 65920 25920 66180
rect 26120 65920 26140 66180
rect 25900 65900 26140 65920
rect 26740 66180 26980 66200
rect 26740 65920 26760 66180
rect 26960 65920 26980 66180
rect 26740 65900 26980 65920
rect 27540 66180 27780 66200
rect 27540 65920 27560 66180
rect 27760 65920 27780 66180
rect 27540 65900 27780 65920
rect 37280 66180 37520 66200
rect 37280 65920 37300 66180
rect 37500 65920 37520 66180
rect 37280 65900 37520 65920
rect 37980 66180 38220 66200
rect 37980 65920 38000 66180
rect 38200 65920 38220 66180
rect 37980 65900 38220 65920
rect 38700 66180 38940 66200
rect 38700 65920 38720 66180
rect 38920 65920 38940 66180
rect 38700 65900 38940 65920
rect 39540 66180 39780 66200
rect 39540 65920 39560 66180
rect 39760 65920 39780 66180
rect 39540 65900 39780 65920
rect 40340 66180 40580 66200
rect 40340 65920 40360 66180
rect 40560 65920 40580 66180
rect 40340 65900 40580 65920
rect 45320 66180 45560 66200
rect 45320 65920 45340 66180
rect 45540 65920 45560 66180
rect 45320 65900 45560 65920
rect 46160 66180 46400 66200
rect 46160 65920 46180 66180
rect 46380 65920 46400 66180
rect 46160 65900 46400 65920
rect 46840 66180 47080 66200
rect 46840 65920 46860 66180
rect 47060 65920 47080 66180
rect 46840 65900 47080 65920
rect 48700 66180 48940 66200
rect 48700 65920 48720 66180
rect 48920 65920 48940 66180
rect 48700 65900 48940 65920
rect 49520 66180 49760 66200
rect 49520 65920 49540 66180
rect 49740 65920 49760 66180
rect 49520 65900 49760 65920
rect 50160 66180 50400 66200
rect 50160 65920 50180 66180
rect 50380 65920 50400 66180
rect 50160 65900 50400 65920
rect 51900 66190 52080 66200
rect 51900 65920 51910 66190
rect 52070 65920 52080 66190
rect 51900 65910 52080 65920
rect 56520 66180 56760 66200
rect 56520 65920 56540 66180
rect 56740 65920 56760 66180
rect 56520 65900 56760 65920
rect 57360 66180 57600 66200
rect 57360 65920 57380 66180
rect 57580 65920 57600 66180
rect 57360 65900 57600 65920
rect 58040 66180 58280 66200
rect 58040 65920 58060 66180
rect 58260 65920 58280 66180
rect 58040 65900 58280 65920
rect 59900 66180 60140 66200
rect 59900 65920 59920 66180
rect 60120 65920 60140 66180
rect 59900 65900 60140 65920
rect 60720 66180 60960 66200
rect 60720 65920 60740 66180
rect 60940 65920 60960 66180
rect 60720 65900 60960 65920
rect 61360 66180 61600 66200
rect 61360 65920 61380 66180
rect 61580 65920 61600 66180
rect 61360 65900 61600 65920
rect 63100 66190 63280 66200
rect 63100 65920 63110 66190
rect 63270 65920 63280 66190
rect 64800 66000 71700 66200
rect 63100 65910 63280 65920
rect 71300 65000 71700 66000
rect 64800 64800 71700 65000
rect 71300 59000 71700 64800
rect 71300 58600 88000 59000
rect 72200 56900 72400 58600
rect 69200 56700 72400 56900
rect 69200 56080 69400 56700
rect 69200 55820 69220 56080
rect 69380 55820 69400 56080
rect 69200 55800 69400 55820
rect 72200 56080 72400 56700
rect 72200 55820 72220 56080
rect 72380 55820 72400 56080
rect 72200 55800 72400 55820
rect 74700 56080 74900 58600
rect 74700 55820 74720 56080
rect 74880 55820 74900 56080
rect 74700 55800 74900 55820
rect 80500 56080 80700 58600
rect 80500 55820 80520 56080
rect 80680 55820 80700 56080
rect 80500 55800 80700 55820
rect 83400 56080 83600 58600
rect 83400 55820 83420 56080
rect 83580 55820 83600 56080
rect 83400 55800 83600 55820
rect 85900 56080 86100 58600
rect 85900 55820 85920 56080
rect 86080 55820 86100 56080
rect 85900 55800 86100 55820
rect 87500 56080 87700 58600
rect 87500 55820 87520 56080
rect 87680 55820 87700 56080
rect 87500 55800 87700 55820
rect 68920 54990 69160 55000
rect 68920 54710 68930 54990
rect 69150 54710 69160 54990
rect 68920 54700 69160 54710
rect 71780 54990 72000 55000
rect 71780 54710 71790 54990
rect 71990 54710 72000 54990
rect 74300 54990 74400 55000
rect 74300 54770 74310 54990
rect 74390 54770 74400 54990
rect 74300 54760 74400 54770
rect 80210 54990 80430 55000
rect 71780 54700 72000 54710
rect 80210 54710 80220 54990
rect 80420 54710 80430 54990
rect 80210 54700 80430 54710
rect 82960 54990 83180 55000
rect 82960 54710 82970 54990
rect 83170 54710 83180 54990
rect 85500 54990 85600 55000
rect 85500 54770 85510 54990
rect 85590 54770 85600 54990
rect 85500 54760 85600 54770
rect 87100 54990 87200 55000
rect 87100 54770 87110 54990
rect 87190 54770 87200 54990
rect 87100 54760 87200 54770
rect 82960 54700 83180 54710
rect 68920 48890 69160 48900
rect 68920 48610 68930 48890
rect 69150 48610 69160 48890
rect 68920 48600 69160 48610
rect 71780 48890 72020 48900
rect 71780 48610 71790 48890
rect 72010 48610 72020 48890
rect 80210 48890 80440 48900
rect 71780 48600 72020 48610
rect 74300 48830 74400 48840
rect 74300 48610 74310 48830
rect 74390 48610 74400 48830
rect 74300 48600 74400 48610
rect 80210 48610 80220 48890
rect 80430 48610 80440 48890
rect 80210 48600 80440 48610
rect 82990 48890 83210 48900
rect 82990 48610 83000 48890
rect 83200 48610 83210 48890
rect 82990 48600 83210 48610
rect 85500 48870 85600 48880
rect 85500 48610 85510 48870
rect 85590 48610 85600 48870
rect 85500 48600 85600 48610
rect 87100 48870 87200 48880
rect 87100 48610 87110 48870
rect 87190 48610 87200 48870
rect 87100 48600 87200 48610
rect 72200 47780 72400 47820
rect 69200 47680 69400 47700
rect 69200 47320 69220 47680
rect 69380 47320 69400 47680
rect 69200 46800 69400 47320
rect 72200 47420 72220 47780
rect 72380 47420 72400 47780
rect 72200 46800 72400 47420
rect 69200 46600 72400 46800
rect 72200 44700 72400 46600
rect 74700 47780 74900 47820
rect 74700 47420 74720 47780
rect 74880 47420 74900 47780
rect 83400 47780 83600 47800
rect 74700 44700 74900 47420
rect 80600 47680 80800 47700
rect 80600 47320 80620 47680
rect 80780 47320 80800 47680
rect 80600 44700 80800 47320
rect 83400 47420 83420 47780
rect 83580 47420 83600 47780
rect 83400 44700 83600 47420
rect 86000 47780 86200 47800
rect 86000 47420 86020 47780
rect 86180 47420 86200 47780
rect 86000 44700 86200 47420
rect 87600 47780 87800 47800
rect 87600 47420 87620 47780
rect 87780 47420 87800 47780
rect 87600 44700 87800 47420
rect 71500 44300 88200 44700
rect 71500 38500 71900 44300
rect 64880 38490 71900 38500
rect 64880 38310 65430 38490
rect 65590 38310 66670 38490
rect 66830 38310 67910 38490
rect 68070 38310 69150 38490
rect 69310 38310 70390 38490
rect 70550 38310 71900 38490
rect 64880 38300 71900 38310
rect -13820 37680 -13540 37700
rect -13820 37420 -13800 37680
rect -13560 37420 -13540 37680
rect -13820 37400 -13540 37420
rect -13120 37680 -12840 37700
rect -13120 37420 -13100 37680
rect -12860 37420 -12840 37680
rect -13120 37400 -12840 37420
rect -12440 37680 -12160 37700
rect -12440 37420 -12420 37680
rect -12180 37420 -12160 37680
rect -12440 37400 -12160 37420
rect -11580 37680 -11300 37700
rect -11580 37420 -11560 37680
rect -11320 37420 -11300 37680
rect -11580 37400 -11300 37420
rect -10800 37680 -10520 37700
rect -10800 37420 -10780 37680
rect -10540 37420 -10520 37680
rect -10800 37400 -10520 37420
rect -1020 37680 -740 37700
rect -1020 37420 -1000 37680
rect -760 37420 -740 37680
rect -1020 37400 -740 37420
rect -380 37680 -100 37700
rect -380 37420 -360 37680
rect -120 37420 -100 37680
rect -380 37400 -100 37420
rect 360 37680 640 37700
rect 360 37420 380 37680
rect 620 37420 640 37680
rect 360 37400 640 37420
rect 1220 37680 1500 37700
rect 1220 37420 1240 37680
rect 1480 37420 1500 37680
rect 1220 37400 1500 37420
rect 2000 37680 2280 37700
rect 2000 37420 2020 37680
rect 2260 37420 2280 37680
rect 2000 37400 2280 37420
rect 24480 37680 24820 37700
rect 24480 37420 24500 37680
rect 24800 37420 24820 37680
rect 24480 37400 24820 37420
rect 25120 37680 25460 37700
rect 25120 37420 25140 37680
rect 25440 37420 25460 37680
rect 25120 37400 25460 37420
rect 25800 37680 26140 37700
rect 25800 37420 25820 37680
rect 26120 37420 26140 37680
rect 25800 37400 26140 37420
rect 26640 37680 26980 37700
rect 26640 37420 26660 37680
rect 26960 37420 26980 37680
rect 26640 37400 26980 37420
rect 27440 37680 27780 37700
rect 27440 37420 27460 37680
rect 27760 37420 27780 37680
rect 27440 37400 27780 37420
rect 37280 37680 37620 37700
rect 37280 37420 37300 37680
rect 37600 37420 37620 37680
rect 37280 37400 37620 37420
rect 37940 37680 38280 37700
rect 37940 37420 37960 37680
rect 38260 37420 38280 37680
rect 37940 37400 38280 37420
rect 38600 37680 38940 37700
rect 38600 37420 38620 37680
rect 38920 37420 38940 37680
rect 38600 37400 38940 37420
rect 39420 37680 39760 37700
rect 39420 37420 39440 37680
rect 39740 37420 39760 37680
rect 39420 37400 39760 37420
rect 40240 37680 40580 37700
rect 40240 37420 40260 37680
rect 40560 37420 40580 37680
rect 40240 37400 40580 37420
rect 45320 37680 45600 37700
rect 45320 37420 45340 37680
rect 45580 37420 45600 37680
rect 45320 37400 45600 37420
rect 46160 37680 46440 37700
rect 46160 37420 46180 37680
rect 46420 37420 46440 37680
rect 46160 37400 46440 37420
rect 46800 37680 47080 37700
rect 46800 37420 46820 37680
rect 47060 37420 47080 37680
rect 46800 37400 47080 37420
rect 48700 37680 49020 37700
rect 48700 37420 48720 37680
rect 49000 37420 49020 37680
rect 48700 37400 49020 37420
rect 49520 37680 49840 37700
rect 49520 37420 49540 37680
rect 49820 37420 49840 37680
rect 49520 37400 49840 37420
rect 50080 37680 50400 37700
rect 50080 37420 50100 37680
rect 50380 37420 50400 37680
rect 50080 37400 50400 37420
rect 51900 37680 52080 37700
rect 51900 37420 51920 37680
rect 52060 37420 52080 37680
rect 51900 37400 52080 37420
rect 56520 37680 56800 37700
rect 56520 37420 56540 37680
rect 56780 37420 56800 37680
rect 56520 37400 56800 37420
rect 57360 37680 57600 37700
rect 57360 37420 57380 37680
rect 57580 37420 57600 37680
rect 57360 37400 57600 37420
rect 58040 37680 58280 37700
rect 58040 37420 58060 37680
rect 58260 37420 58280 37680
rect 58040 37400 58280 37420
rect 59900 37680 60120 37700
rect 59900 37420 59920 37680
rect 60100 37420 60120 37680
rect 59900 37400 60120 37420
rect 60720 37680 60940 37700
rect 60720 37420 60740 37680
rect 60920 37420 60940 37680
rect 60720 37400 60940 37420
rect 61380 37680 61600 37700
rect 61380 37420 61400 37680
rect 61580 37420 61600 37680
rect 61380 37400 61600 37420
rect 63100 37640 63280 37660
rect 63100 37420 63120 37640
rect 63260 37420 63280 37640
rect 71500 37500 71900 38300
rect 63100 37400 63280 37420
rect 64880 37490 71900 37500
rect 64880 37310 65430 37490
rect 65590 37310 66670 37490
rect 66830 37310 67910 37490
rect 68070 37310 69150 37490
rect 69310 37310 70390 37490
rect 70550 37310 71900 37490
rect 64880 37300 71900 37310
rect 52200 36580 52400 36600
rect -13400 36180 -13200 36200
rect -13400 35820 -13380 36180
rect -13220 35820 -13200 36180
rect -13400 33400 -13200 35820
rect -600 36180 -400 36200
rect -600 35820 -580 36180
rect -420 35820 -400 36180
rect -600 33400 -400 35820
rect 24800 36180 25000 36200
rect 24800 35820 24820 36180
rect 24980 35820 25000 36180
rect 24800 33400 25000 35820
rect 27100 33400 27300 36300
rect 37600 36180 37800 36200
rect 37600 35820 37620 36180
rect 37780 35820 37800 36180
rect 37600 33400 37800 35820
rect 39900 33400 40100 36300
rect 45400 33400 45600 36300
rect 46800 36180 47000 36200
rect 46800 35820 46820 36180
rect 46980 35820 47000 36180
rect 46800 33400 47000 35820
rect 48700 33400 48900 36300
rect 50200 36180 50400 36200
rect 50200 35820 50220 36180
rect 50380 35820 50400 36180
rect 50200 33400 50400 35820
rect 51500 33400 51700 36500
rect 52200 36220 52220 36580
rect 52380 36220 52400 36580
rect 52200 33400 52400 36220
rect 56600 33400 56800 36300
rect 58000 36180 58200 36200
rect 58000 35820 58020 36180
rect 58180 35820 58200 36180
rect 58000 33400 58200 35820
rect 60000 33400 60200 36300
rect 61400 36180 61600 36200
rect 61400 35820 61420 36180
rect 61580 35820 61600 36180
rect 61400 33400 61600 35820
rect 62600 33400 62800 36600
rect 63400 36580 63600 36600
rect 63400 36220 63420 36580
rect 63580 36220 63600 36580
rect 63400 33400 63600 36220
rect 71500 33400 71900 37300
rect -13400 33000 71900 33400
<< via3 >>
rect -13800 65920 -13600 66180
rect -13120 65920 -12920 66180
rect -12380 65920 -12180 66180
rect -11540 65920 -11340 66180
rect -10740 65920 -10540 66180
rect -1000 65920 -820 66180
rect -300 65920 -120 66180
rect 440 65920 620 66180
rect 1220 65920 1400 66180
rect 2060 65920 2240 66180
rect 24500 65920 24700 66180
rect 25200 65920 25400 66180
rect 25920 65920 26120 66180
rect 26760 65920 26960 66180
rect 27560 65920 27760 66180
rect 37300 65920 37500 66180
rect 38000 65920 38200 66180
rect 38720 65920 38920 66180
rect 39560 65920 39760 66180
rect 40360 65920 40560 66180
rect 45340 65920 45540 66180
rect 46180 65920 46380 66180
rect 46860 65920 47060 66180
rect 48720 65920 48920 66180
rect 49540 65920 49740 66180
rect 50180 65920 50380 66180
rect 51910 65920 52070 66190
rect 56540 65920 56740 66180
rect 57380 65920 57580 66180
rect 58060 65920 58260 66180
rect 59920 65920 60120 66180
rect 60740 65920 60940 66180
rect 61380 65920 61580 66180
rect 63110 65920 63270 66190
rect 68930 54710 69150 54990
rect 71790 54710 71990 54990
rect 74310 54770 74390 54990
rect 80220 54710 80420 54990
rect 82970 54710 83170 54990
rect 85510 54770 85590 54990
rect 87110 54770 87190 54990
rect 68930 48610 69150 48890
rect 71790 48610 72010 48890
rect 74310 48610 74390 48830
rect 80220 48610 80430 48890
rect 83000 48610 83200 48890
rect 85510 48610 85590 48870
rect 87110 48610 87190 48870
rect -13800 37420 -13560 37680
rect -13100 37420 -12860 37680
rect -12420 37420 -12180 37680
rect -11560 37420 -11320 37680
rect -10780 37420 -10540 37680
rect -1000 37420 -760 37680
rect -360 37420 -120 37680
rect 380 37420 620 37680
rect 1240 37420 1480 37680
rect 2020 37420 2260 37680
rect 24500 37420 24800 37680
rect 25140 37420 25440 37680
rect 25820 37420 26120 37680
rect 26660 37420 26960 37680
rect 27460 37420 27760 37680
rect 37300 37420 37600 37680
rect 37960 37420 38260 37680
rect 38620 37420 38920 37680
rect 39440 37420 39740 37680
rect 40260 37420 40560 37680
rect 45340 37420 45580 37680
rect 46180 37420 46420 37680
rect 46820 37420 47060 37680
rect 48720 37420 49000 37680
rect 49540 37420 49820 37680
rect 50100 37420 50380 37680
rect 51920 37420 52060 37680
rect 56540 37420 56780 37680
rect 57380 37420 57580 37680
rect 58060 37420 58260 37680
rect 59920 37420 60100 37680
rect 60740 37420 60920 37680
rect 61400 37420 61580 37680
rect 63120 37420 63260 37640
<< metal4 >>
rect 51900 66190 52080 66200
rect 51900 65920 51910 66190
rect 52070 65920 52080 66190
rect 63100 66190 63280 66200
rect 63100 65920 63110 66190
rect 63270 65920 63280 66190
rect 51900 65910 52080 65920
rect 63100 65910 63280 65920
rect 71500 44300 88200 44700
rect 51900 37680 52080 37700
rect 51900 37420 51920 37680
rect 52060 37420 52080 37680
rect 63100 37640 63280 37660
rect 63100 37420 63120 37640
rect 63260 37420 63280 37640
rect 51900 37400 52080 37420
rect 63100 37400 63280 37420
rect -11100 33400 -10900 36300
rect 1600 33400 1800 36300
rect 27100 33400 27300 36300
rect 39900 33400 40100 36300
rect 45400 33400 45600 36300
rect 48700 33400 48900 36300
rect 51500 33400 51700 36500
rect 56600 33400 56800 36300
rect 60000 33400 60200 36300
rect 62600 33400 62800 36600
rect 71500 33400 71900 44300
rect -13400 33000 71900 33400
use capacitor_array  capacitor_array_0
timestamp 1667870970
transform 1 0 0 0 1 40400
box -35000 -3000 87900 25800
use capacitor_switch2  capacitor_switch2_0
timestamp 1668018737
transform 0 -1 88140 1 0 47570
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_1
timestamp 1668018737
transform 0 -1 72840 1 0 47570
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_2
timestamp 1668018737
transform 0 -1 75290 1 0 47570
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_3
timestamp 1668018737
transform 0 -1 84040 1 0 47570
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_4
timestamp 1668018737
transform 0 -1 86540 1 0 47570
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_5
timestamp 1668018737
transform 0 -1 75340 -1 0 55930
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_6
timestamp 1668018737
transform 0 -1 72840 -1 0 55930
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_7
timestamp 1668018737
transform 0 -1 84040 -1 0 55930
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_8
timestamp 1668018737
transform 0 -1 86540 -1 0 55930
box -300 650 730 1240
use capacitor_switch2  capacitor_switch2_9
timestamp 1668018737
transform 0 -1 88140 -1 0 55930
box -300 650 730 1240
use capacitor_switch4  capacitor_switch4_0
timestamp 1668017310
transform 0 -1 64110 1 0 35900
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_1
timestamp 1668017310
transform 0 -1 81270 1 0 47000
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_2
timestamp 1668017310
transform 0 -1 52960 1 0 35900
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_3
timestamp 1668017310
transform 0 -1 69970 1 0 47000
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_4
timestamp 1668017310
transform 0 -1 69970 -1 0 56500
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_5
timestamp 1668017310
transform 0 -1 81270 -1 0 56500
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_6
timestamp 1668017310
transform 0 -1 64170 -1 0 67700
box 200 530 1300 1570
use capacitor_switch4  capacitor_switch4_7
timestamp 1668017310
transform 0 -1 52960 -1 0 67700
box 200 530 1300 1570
use capacitor_switch8  capacitor_switch8_0
timestamp 1668016891
transform 0 -1 58460 -1 0 68380
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_1
timestamp 1668016891
transform 0 -1 47260 -1 0 68380
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_2
timestamp 1668016891
transform 0 -1 50620 -1 0 68380
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_3
timestamp 1668016891
transform 0 -1 61820 -1 0 68380
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_4
timestamp 1668016891
transform 0 -1 50620 1 0 35220
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_5
timestamp 1668016891
transform 0 -1 47260 1 0 35220
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_6
timestamp 1668016891
transform 0 -1 58460 1 0 35220
box -20 90 1980 2060
use capacitor_switch8  capacitor_switch8_7
timestamp 1668016891
transform 0 -1 61820 1 0 35220
box -20 90 1980 2060
use capacitor_switch16  capacitor_switch16_0
timestamp 1668016263
transform 0 1 -13250 -1 0 68090
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_1
timestamp 1668016263
transform 0 1 37850 -1 0 68090
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_2
timestamp 1668016263
transform 0 1 -450 -1 0 68090
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_3
timestamp 1668016263
transform 0 1 25050 -1 0 68090
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_4
timestamp 1668016263
transform 0 1 -450 1 0 35510
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_5
timestamp 1668016263
transform 0 1 -13250 1 0 35510
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_6
timestamp 1668016263
transform 0 1 25050 1 0 35510
box -300 -650 1730 2810
use capacitor_switch16  capacitor_switch16_7
timestamp 1668016263
transform 0 1 37850 1 0 35510
box -300 -650 1730 2810
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 0 1 65548 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_1
timestamp 1662439860
transform 0 -1 69192 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_2
timestamp 1662439860
transform 0 -1 67952 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_3
timestamp 1662439860
transform 0 -1 66712 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_4
timestamp 1662439860
transform 0 -1 65472 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_5
timestamp 1662439860
transform 0 1 70508 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_6
timestamp 1662439860
transform 0 1 68028 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_7
timestamp 1662439860
transform 0 1 66788 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_8
timestamp 1662439860
transform 0 1 69268 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_9
timestamp 1662439860
transform 0 -1 70432 -1 0 39362
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_10
timestamp 1662439860
transform 0 1 65548 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_11
timestamp 1662439860
transform 0 -1 66712 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_12
timestamp 1662439860
transform 0 -1 65472 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_13
timestamp 1662439860
transform 0 1 66788 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_14
timestamp 1662439860
transform 0 -1 67952 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_15
timestamp 1662439860
transform 0 1 68028 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_16
timestamp 1662439860
transform 0 -1 69192 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_17
timestamp 1662439860
transform 0 1 70508 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_18
timestamp 1662439860
transform 0 1 69268 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  sky130_fd_sc_hd__bufbuf_16_19
timestamp 1662439860
transform 0 -1 70432 1 0 64038
box -38 -48 2430 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 0 -1 66712 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_1
timestamp 1662439860
transform 0 -1 65472 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_2
timestamp 1662439860
transform 0 -1 69192 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_3
timestamp 1662439860
transform 0 -1 67952 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_4
timestamp 1662439860
transform 0 -1 70432 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_5
timestamp 1662439860
transform 0 1 65548 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_6
timestamp 1662439860
transform 0 1 66788 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_7
timestamp 1662439860
transform 0 1 68028 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_8
timestamp 1662439860
transform 0 1 70508 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_9
timestamp 1662439860
transform 0 1 69268 1 0 63578
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_10
timestamp 1662439860
transform 0 -1 67952 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_11
timestamp 1662439860
transform 0 1 66788 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_12
timestamp 1662439860
transform 0 -1 66712 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_13
timestamp 1662439860
transform 0 1 65548 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_14
timestamp 1662439860
transform 0 -1 65472 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_15
timestamp 1662439860
transform 0 1 70508 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_16
timestamp 1662439860
transform 0 -1 70432 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_17
timestamp 1662439860
transform 0 1 69268 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_18
timestamp 1662439860
transform 0 -1 69192 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_19
timestamp 1662439860
transform 0 1 68028 1 0 36688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_20
timestamp 1662439860
transform 0 -1 65472 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_21
timestamp 1662439860
transform 0 -1 66712 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_22
timestamp 1662439860
transform 0 1 65548 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_23
timestamp 1662439860
transform 0 -1 67952 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_24
timestamp 1662439860
transform 0 1 66788 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_25
timestamp 1662439860
transform 0 -1 69192 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_26
timestamp 1662439860
transform 0 1 68028 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_27
timestamp 1662439860
transform 0 -1 70432 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_28
timestamp 1662439860
transform 0 1 69268 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_29
timestamp 1662439860
transform 0 1 70508 -1 0 66712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_30
timestamp 1662439860
transform 0 1 70508 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_31
timestamp 1662439860
transform 0 -1 70432 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_32
timestamp 1662439860
transform 0 1 69268 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_33
timestamp 1662439860
transform 0 -1 69192 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_34
timestamp 1662439860
transform 0 1 68028 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_35
timestamp 1662439860
transform 0 -1 67952 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_36
timestamp 1662439860
transform 0 1 66788 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_37
timestamp 1662439860
transform 0 -1 66712 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_38
timestamp 1662439860
transform 0 -1 65472 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_39
timestamp 1662439860
transform 0 1 65548 -1 0 39822
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 0 1 65548 1 0 39450
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1662439860
transform 0 -1 66712 -1 0 39542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1662439860
transform 0 -1 69192 -1 0 39542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1662439860
transform 0 -1 67952 -1 0 39542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1662439860
transform 0 -1 70432 -1 0 39542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1662439860
transform 0 -1 65472 -1 0 39542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1662439860
transform 0 1 69268 1 0 39450
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1662439860
transform 0 1 66788 1 0 39450
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1662439860
transform 0 1 68028 1 0 39450
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1662439860
transform 0 1 70508 1 0 39450
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1662439860
transform 0 1 65548 -1 0 63950
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1662439860
transform 0 -1 66712 1 0 63858
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1662439860
transform 0 -1 65472 1 0 63858
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1662439860
transform 0 1 66788 -1 0 63950
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1662439860
transform 0 -1 67952 1 0 63858
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1662439860
transform 0 1 68028 -1 0 63950
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1662439860
transform 0 -1 69192 1 0 63858
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1662439860
transform 0 -1 70432 1 0 63858
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1662439860
transform 0 1 69268 -1 0 63950
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1662439860
transform 0 1 70508 -1 0 63950
box -38 -48 130 592
<< labels >>
flabel nwell s 71035 64028 71069 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 64048 71069 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 64038 71069 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 64058 71069 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 64078 71069 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 39288 71069 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 39308 71069 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 39328 71069 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 39318 71069 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 71035 39338 71069 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 64028 69809 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 64028 69905 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 64048 69905 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 64048 69809 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 64068 69849 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 64028 69829 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 64028 69849 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 64048 69849 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 64048 69829 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 63607 69829 63641 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 64068 69829 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 66649 69829 66683 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 64038 69809 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 64038 69905 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 64058 69905 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 64058 69809 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 64078 69849 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 64038 69829 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 64038 69849 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 64058 69849 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 64058 69829 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 64078 69829 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 64078 69809 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 64078 69905 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 64028 68569 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 64028 68665 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 64048 68569 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 64048 68665 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 64068 68609 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 64028 68589 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 64028 68609 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 64048 68609 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 64048 68589 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 63607 68589 63641 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 64068 68589 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 66649 68589 66683 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 64038 68569 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 64038 68665 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 64058 68569 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 64058 68665 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 64078 68609 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 64038 68589 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 64038 68609 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 64058 68609 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 64058 68589 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 64078 68589 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 64078 68569 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 64078 68665 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 64028 67329 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 64028 67425 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 64048 67329 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 64048 67425 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 64068 67369 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 64028 67349 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 64028 67369 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 64048 67369 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 64048 67349 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 63607 67349 63641 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 64068 67349 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 66649 67349 66683 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 64038 67329 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 64038 67425 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 64058 67329 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 64058 67425 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 64078 67369 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 64038 67349 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 64038 67369 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 64058 67369 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 64058 67349 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 64078 67349 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 64078 67329 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 64078 67425 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 64028 66089 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 64028 66185 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 64048 66089 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 64048 66185 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 64068 66129 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 64028 66109 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 64028 66129 64062 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 64048 66129 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 64048 66109 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 63607 66109 63641 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 64068 66109 64102 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 66649 66109 66683 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 64038 66089 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 64038 66185 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 64058 66089 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 64058 66185 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 64078 66129 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 64038 66109 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 64038 66129 64072 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 64058 66129 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 64058 66109 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 64078 66109 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 64078 66089 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 64078 66185 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 64911 64048 64945 64082 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 64911 64058 64945 64092 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 64911 64078 64945 64112 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 39288 69905 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 39288 69809 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39288 69829 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39308 69829 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 39308 69849 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 39328 69849 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39328 69829 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 39288 69849 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 39308 69809 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 39308 69905 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 39328 69905 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 39328 69809 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 36717 69829 36751 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39298 69829 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39759 69829 39793 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39318 69829 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 39318 69849 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 39338 69849 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69795 39338 69829 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69815 39298 69849 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 39318 69809 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 39318 69905 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69871 39338 69905 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 69775 39338 69809 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 39288 68665 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 39288 68569 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39288 68589 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39308 68589 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 39308 68609 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 39328 68609 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39328 68589 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 39288 68609 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 39308 68665 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 39308 68569 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 39328 68665 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 39328 68569 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 36717 68589 36751 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39298 68589 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39759 68589 39793 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39318 68589 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 39318 68609 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 39338 68609 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68555 39338 68589 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68575 39298 68609 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 39318 68665 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 39318 68569 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68631 39338 68665 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 68535 39338 68569 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 39288 67425 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 39288 67329 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39288 67349 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39308 67349 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 39308 67369 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 39328 67369 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39328 67349 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 39288 67369 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 39308 67425 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 39308 67329 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 39328 67425 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 39328 67329 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 36717 67349 36751 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39298 67349 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39759 67349 39793 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39318 67349 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 39318 67369 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 39338 67369 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67315 39338 67349 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67335 39298 67369 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 39318 67425 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 39318 67329 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67391 39338 67425 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 67295 39338 67329 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 39288 66185 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 39288 66089 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39288 66109 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39308 66109 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 39308 66129 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 39328 66129 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39328 66109 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 39288 66129 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 39308 66185 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 39308 66089 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 39328 66185 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 39328 66089 39362 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 36717 66109 36751 0 FreeSans 200 270 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39298 66109 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39759 66109 39793 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39318 66109 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 39318 66129 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 39338 66129 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66075 39338 66109 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66095 39298 66129 39332 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 39318 66185 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 39318 66089 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66151 39338 66185 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 66055 39338 66089 39372 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 64911 39318 64945 39352 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 64911 39308 64945 39342 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 64911 39288 64945 39322 0 FreeSans 200 90 0 0 VPB
port 4 nsew power bidirectional
<< end >>
