magic
tech sky130A
magscale 1 2
timestamp 1666651042
<< nmos >>
rect -15 -91 15 91
<< ndiff >>
rect -73 79 -15 91
rect -73 -79 -61 79
rect -27 -79 -15 79
rect -73 -91 -15 -79
rect 15 79 73 91
rect 15 -79 27 79
rect 61 -79 73 79
rect 15 -91 73 -79
<< ndiffc >>
rect -61 -79 -27 79
rect 27 -79 61 79
<< poly >>
rect -15 91 15 117
rect -15 -117 15 -91
<< locali >>
rect -61 79 -27 95
rect -61 -95 -27 -79
rect 27 79 61 95
rect 27 -95 61 -79
<< viali >>
rect -61 -79 -27 79
rect 27 -79 61 79
<< metal1 >>
rect -67 79 -21 91
rect -67 -79 -61 79
rect -27 -79 -21 79
rect -67 -91 -21 -79
rect 21 79 67 91
rect 21 -79 27 79
rect 61 -79 67 79
rect 21 -91 67 -79
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
