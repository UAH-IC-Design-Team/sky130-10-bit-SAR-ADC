magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< metal3 >>
rect -350 288562 349 288590
rect -350 284208 265 288562
rect 329 284208 349 288562
rect -350 284180 349 284208
rect -350 284052 349 284080
rect -350 279698 265 284052
rect 329 279698 349 284052
rect -350 279670 349 279698
rect -350 279542 349 279570
rect -350 275188 265 279542
rect 329 275188 349 279542
rect -350 275160 349 275188
rect -350 275032 349 275060
rect -350 270678 265 275032
rect 329 270678 349 275032
rect -350 270650 349 270678
rect -350 270522 349 270550
rect -350 266168 265 270522
rect 329 266168 349 270522
rect -350 266140 349 266168
rect -350 266012 349 266040
rect -350 261658 265 266012
rect 329 261658 349 266012
rect -350 261630 349 261658
rect -350 261502 349 261530
rect -350 257148 265 261502
rect 329 257148 349 261502
rect -350 257120 349 257148
rect -350 256992 349 257020
rect -350 252638 265 256992
rect 329 252638 349 256992
rect -350 252610 349 252638
rect -350 252482 349 252510
rect -350 248128 265 252482
rect 329 248128 349 252482
rect -350 248100 349 248128
rect -350 247972 349 248000
rect -350 243618 265 247972
rect 329 243618 349 247972
rect -350 243590 349 243618
rect -350 243462 349 243490
rect -350 239108 265 243462
rect 329 239108 349 243462
rect -350 239080 349 239108
rect -350 238952 349 238980
rect -350 234598 265 238952
rect 329 234598 349 238952
rect -350 234570 349 234598
rect -350 234442 349 234470
rect -350 230088 265 234442
rect 329 230088 349 234442
rect -350 230060 349 230088
rect -350 229932 349 229960
rect -350 225578 265 229932
rect 329 225578 349 229932
rect -350 225550 349 225578
rect -350 225422 349 225450
rect -350 221068 265 225422
rect 329 221068 349 225422
rect -350 221040 349 221068
rect -350 220912 349 220940
rect -350 216558 265 220912
rect 329 216558 349 220912
rect -350 216530 349 216558
rect -350 216402 349 216430
rect -350 212048 265 216402
rect 329 212048 349 216402
rect -350 212020 349 212048
rect -350 211892 349 211920
rect -350 207538 265 211892
rect 329 207538 349 211892
rect -350 207510 349 207538
rect -350 207382 349 207410
rect -350 203028 265 207382
rect 329 203028 349 207382
rect -350 203000 349 203028
rect -350 202872 349 202900
rect -350 198518 265 202872
rect 329 198518 349 202872
rect -350 198490 349 198518
rect -350 198362 349 198390
rect -350 194008 265 198362
rect 329 194008 349 198362
rect -350 193980 349 194008
rect -350 193852 349 193880
rect -350 189498 265 193852
rect 329 189498 349 193852
rect -350 189470 349 189498
rect -350 189342 349 189370
rect -350 184988 265 189342
rect 329 184988 349 189342
rect -350 184960 349 184988
rect -350 184832 349 184860
rect -350 180478 265 184832
rect 329 180478 349 184832
rect -350 180450 349 180478
rect -350 180322 349 180350
rect -350 175968 265 180322
rect 329 175968 349 180322
rect -350 175940 349 175968
rect -350 175812 349 175840
rect -350 171458 265 175812
rect 329 171458 349 175812
rect -350 171430 349 171458
rect -350 171302 349 171330
rect -350 166948 265 171302
rect 329 166948 349 171302
rect -350 166920 349 166948
rect -350 166792 349 166820
rect -350 162438 265 166792
rect 329 162438 349 166792
rect -350 162410 349 162438
rect -350 162282 349 162310
rect -350 157928 265 162282
rect 329 157928 349 162282
rect -350 157900 349 157928
rect -350 157772 349 157800
rect -350 153418 265 157772
rect 329 153418 349 157772
rect -350 153390 349 153418
rect -350 153262 349 153290
rect -350 148908 265 153262
rect 329 148908 349 153262
rect -350 148880 349 148908
rect -350 148752 349 148780
rect -350 144398 265 148752
rect 329 144398 349 148752
rect -350 144370 349 144398
rect -350 144242 349 144270
rect -350 139888 265 144242
rect 329 139888 349 144242
rect -350 139860 349 139888
rect -350 139732 349 139760
rect -350 135378 265 139732
rect 329 135378 349 139732
rect -350 135350 349 135378
rect -350 135222 349 135250
rect -350 130868 265 135222
rect 329 130868 349 135222
rect -350 130840 349 130868
rect -350 130712 349 130740
rect -350 126358 265 130712
rect 329 126358 349 130712
rect -350 126330 349 126358
rect -350 126202 349 126230
rect -350 121848 265 126202
rect 329 121848 349 126202
rect -350 121820 349 121848
rect -350 121692 349 121720
rect -350 117338 265 121692
rect 329 117338 349 121692
rect -350 117310 349 117338
rect -350 117182 349 117210
rect -350 112828 265 117182
rect 329 112828 349 117182
rect -350 112800 349 112828
rect -350 112672 349 112700
rect -350 108318 265 112672
rect 329 108318 349 112672
rect -350 108290 349 108318
rect -350 108162 349 108190
rect -350 103808 265 108162
rect 329 103808 349 108162
rect -350 103780 349 103808
rect -350 103652 349 103680
rect -350 99298 265 103652
rect 329 99298 349 103652
rect -350 99270 349 99298
rect -350 99142 349 99170
rect -350 94788 265 99142
rect 329 94788 349 99142
rect -350 94760 349 94788
rect -350 94632 349 94660
rect -350 90278 265 94632
rect 329 90278 349 94632
rect -350 90250 349 90278
rect -350 90122 349 90150
rect -350 85768 265 90122
rect 329 85768 349 90122
rect -350 85740 349 85768
rect -350 85612 349 85640
rect -350 81258 265 85612
rect 329 81258 349 85612
rect -350 81230 349 81258
rect -350 81102 349 81130
rect -350 76748 265 81102
rect 329 76748 349 81102
rect -350 76720 349 76748
rect -350 76592 349 76620
rect -350 72238 265 76592
rect 329 72238 349 76592
rect -350 72210 349 72238
rect -350 72082 349 72110
rect -350 67728 265 72082
rect 329 67728 349 72082
rect -350 67700 349 67728
rect -350 67572 349 67600
rect -350 63218 265 67572
rect 329 63218 349 67572
rect -350 63190 349 63218
rect -350 63062 349 63090
rect -350 58708 265 63062
rect 329 58708 349 63062
rect -350 58680 349 58708
rect -350 58552 349 58580
rect -350 54198 265 58552
rect 329 54198 349 58552
rect -350 54170 349 54198
rect -350 54042 349 54070
rect -350 49688 265 54042
rect 329 49688 349 54042
rect -350 49660 349 49688
rect -350 49532 349 49560
rect -350 45178 265 49532
rect 329 45178 349 49532
rect -350 45150 349 45178
rect -350 45022 349 45050
rect -350 40668 265 45022
rect 329 40668 349 45022
rect -350 40640 349 40668
rect -350 40512 349 40540
rect -350 36158 265 40512
rect 329 36158 349 40512
rect -350 36130 349 36158
rect -350 36002 349 36030
rect -350 31648 265 36002
rect 329 31648 349 36002
rect -350 31620 349 31648
rect -350 31492 349 31520
rect -350 27138 265 31492
rect 329 27138 349 31492
rect -350 27110 349 27138
rect -350 26982 349 27010
rect -350 22628 265 26982
rect 329 22628 349 26982
rect -350 22600 349 22628
rect -350 22472 349 22500
rect -350 18118 265 22472
rect 329 18118 349 22472
rect -350 18090 349 18118
rect -350 17962 349 17990
rect -350 13608 265 17962
rect 329 13608 349 17962
rect -350 13580 349 13608
rect -350 13452 349 13480
rect -350 9098 265 13452
rect 329 9098 349 13452
rect -350 9070 349 9098
rect -350 8942 349 8970
rect -350 4588 265 8942
rect 329 4588 349 8942
rect -350 4560 349 4588
rect -350 4432 349 4460
rect -350 78 265 4432
rect 329 78 349 4432
rect -350 50 349 78
rect -350 -78 349 -50
rect -350 -4432 265 -78
rect 329 -4432 349 -78
rect -350 -4460 349 -4432
rect -350 -4588 349 -4560
rect -350 -8942 265 -4588
rect 329 -8942 349 -4588
rect -350 -8970 349 -8942
rect -350 -9098 349 -9070
rect -350 -13452 265 -9098
rect 329 -13452 349 -9098
rect -350 -13480 349 -13452
rect -350 -13608 349 -13580
rect -350 -17962 265 -13608
rect 329 -17962 349 -13608
rect -350 -17990 349 -17962
rect -350 -18118 349 -18090
rect -350 -22472 265 -18118
rect 329 -22472 349 -18118
rect -350 -22500 349 -22472
rect -350 -22628 349 -22600
rect -350 -26982 265 -22628
rect 329 -26982 349 -22628
rect -350 -27010 349 -26982
rect -350 -27138 349 -27110
rect -350 -31492 265 -27138
rect 329 -31492 349 -27138
rect -350 -31520 349 -31492
rect -350 -31648 349 -31620
rect -350 -36002 265 -31648
rect 329 -36002 349 -31648
rect -350 -36030 349 -36002
rect -350 -36158 349 -36130
rect -350 -40512 265 -36158
rect 329 -40512 349 -36158
rect -350 -40540 349 -40512
rect -350 -40668 349 -40640
rect -350 -45022 265 -40668
rect 329 -45022 349 -40668
rect -350 -45050 349 -45022
rect -350 -45178 349 -45150
rect -350 -49532 265 -45178
rect 329 -49532 349 -45178
rect -350 -49560 349 -49532
rect -350 -49688 349 -49660
rect -350 -54042 265 -49688
rect 329 -54042 349 -49688
rect -350 -54070 349 -54042
rect -350 -54198 349 -54170
rect -350 -58552 265 -54198
rect 329 -58552 349 -54198
rect -350 -58580 349 -58552
rect -350 -58708 349 -58680
rect -350 -63062 265 -58708
rect 329 -63062 349 -58708
rect -350 -63090 349 -63062
rect -350 -63218 349 -63190
rect -350 -67572 265 -63218
rect 329 -67572 349 -63218
rect -350 -67600 349 -67572
rect -350 -67728 349 -67700
rect -350 -72082 265 -67728
rect 329 -72082 349 -67728
rect -350 -72110 349 -72082
rect -350 -72238 349 -72210
rect -350 -76592 265 -72238
rect 329 -76592 349 -72238
rect -350 -76620 349 -76592
rect -350 -76748 349 -76720
rect -350 -81102 265 -76748
rect 329 -81102 349 -76748
rect -350 -81130 349 -81102
rect -350 -81258 349 -81230
rect -350 -85612 265 -81258
rect 329 -85612 349 -81258
rect -350 -85640 349 -85612
rect -350 -85768 349 -85740
rect -350 -90122 265 -85768
rect 329 -90122 349 -85768
rect -350 -90150 349 -90122
rect -350 -90278 349 -90250
rect -350 -94632 265 -90278
rect 329 -94632 349 -90278
rect -350 -94660 349 -94632
rect -350 -94788 349 -94760
rect -350 -99142 265 -94788
rect 329 -99142 349 -94788
rect -350 -99170 349 -99142
rect -350 -99298 349 -99270
rect -350 -103652 265 -99298
rect 329 -103652 349 -99298
rect -350 -103680 349 -103652
rect -350 -103808 349 -103780
rect -350 -108162 265 -103808
rect 329 -108162 349 -103808
rect -350 -108190 349 -108162
rect -350 -108318 349 -108290
rect -350 -112672 265 -108318
rect 329 -112672 349 -108318
rect -350 -112700 349 -112672
rect -350 -112828 349 -112800
rect -350 -117182 265 -112828
rect 329 -117182 349 -112828
rect -350 -117210 349 -117182
rect -350 -117338 349 -117310
rect -350 -121692 265 -117338
rect 329 -121692 349 -117338
rect -350 -121720 349 -121692
rect -350 -121848 349 -121820
rect -350 -126202 265 -121848
rect 329 -126202 349 -121848
rect -350 -126230 349 -126202
rect -350 -126358 349 -126330
rect -350 -130712 265 -126358
rect 329 -130712 349 -126358
rect -350 -130740 349 -130712
rect -350 -130868 349 -130840
rect -350 -135222 265 -130868
rect 329 -135222 349 -130868
rect -350 -135250 349 -135222
rect -350 -135378 349 -135350
rect -350 -139732 265 -135378
rect 329 -139732 349 -135378
rect -350 -139760 349 -139732
rect -350 -139888 349 -139860
rect -350 -144242 265 -139888
rect 329 -144242 349 -139888
rect -350 -144270 349 -144242
rect -350 -144398 349 -144370
rect -350 -148752 265 -144398
rect 329 -148752 349 -144398
rect -350 -148780 349 -148752
rect -350 -148908 349 -148880
rect -350 -153262 265 -148908
rect 329 -153262 349 -148908
rect -350 -153290 349 -153262
rect -350 -153418 349 -153390
rect -350 -157772 265 -153418
rect 329 -157772 349 -153418
rect -350 -157800 349 -157772
rect -350 -157928 349 -157900
rect -350 -162282 265 -157928
rect 329 -162282 349 -157928
rect -350 -162310 349 -162282
rect -350 -162438 349 -162410
rect -350 -166792 265 -162438
rect 329 -166792 349 -162438
rect -350 -166820 349 -166792
rect -350 -166948 349 -166920
rect -350 -171302 265 -166948
rect 329 -171302 349 -166948
rect -350 -171330 349 -171302
rect -350 -171458 349 -171430
rect -350 -175812 265 -171458
rect 329 -175812 349 -171458
rect -350 -175840 349 -175812
rect -350 -175968 349 -175940
rect -350 -180322 265 -175968
rect 329 -180322 349 -175968
rect -350 -180350 349 -180322
rect -350 -180478 349 -180450
rect -350 -184832 265 -180478
rect 329 -184832 349 -180478
rect -350 -184860 349 -184832
rect -350 -184988 349 -184960
rect -350 -189342 265 -184988
rect 329 -189342 349 -184988
rect -350 -189370 349 -189342
rect -350 -189498 349 -189470
rect -350 -193852 265 -189498
rect 329 -193852 349 -189498
rect -350 -193880 349 -193852
rect -350 -194008 349 -193980
rect -350 -198362 265 -194008
rect 329 -198362 349 -194008
rect -350 -198390 349 -198362
rect -350 -198518 349 -198490
rect -350 -202872 265 -198518
rect 329 -202872 349 -198518
rect -350 -202900 349 -202872
rect -350 -203028 349 -203000
rect -350 -207382 265 -203028
rect 329 -207382 349 -203028
rect -350 -207410 349 -207382
rect -350 -207538 349 -207510
rect -350 -211892 265 -207538
rect 329 -211892 349 -207538
rect -350 -211920 349 -211892
rect -350 -212048 349 -212020
rect -350 -216402 265 -212048
rect 329 -216402 349 -212048
rect -350 -216430 349 -216402
rect -350 -216558 349 -216530
rect -350 -220912 265 -216558
rect 329 -220912 349 -216558
rect -350 -220940 349 -220912
rect -350 -221068 349 -221040
rect -350 -225422 265 -221068
rect 329 -225422 349 -221068
rect -350 -225450 349 -225422
rect -350 -225578 349 -225550
rect -350 -229932 265 -225578
rect 329 -229932 349 -225578
rect -350 -229960 349 -229932
rect -350 -230088 349 -230060
rect -350 -234442 265 -230088
rect 329 -234442 349 -230088
rect -350 -234470 349 -234442
rect -350 -234598 349 -234570
rect -350 -238952 265 -234598
rect 329 -238952 349 -234598
rect -350 -238980 349 -238952
rect -350 -239108 349 -239080
rect -350 -243462 265 -239108
rect 329 -243462 349 -239108
rect -350 -243490 349 -243462
rect -350 -243618 349 -243590
rect -350 -247972 265 -243618
rect 329 -247972 349 -243618
rect -350 -248000 349 -247972
rect -350 -248128 349 -248100
rect -350 -252482 265 -248128
rect 329 -252482 349 -248128
rect -350 -252510 349 -252482
rect -350 -252638 349 -252610
rect -350 -256992 265 -252638
rect 329 -256992 349 -252638
rect -350 -257020 349 -256992
rect -350 -257148 349 -257120
rect -350 -261502 265 -257148
rect 329 -261502 349 -257148
rect -350 -261530 349 -261502
rect -350 -261658 349 -261630
rect -350 -266012 265 -261658
rect 329 -266012 349 -261658
rect -350 -266040 349 -266012
rect -350 -266168 349 -266140
rect -350 -270522 265 -266168
rect 329 -270522 349 -266168
rect -350 -270550 349 -270522
rect -350 -270678 349 -270650
rect -350 -275032 265 -270678
rect 329 -275032 349 -270678
rect -350 -275060 349 -275032
rect -350 -275188 349 -275160
rect -350 -279542 265 -275188
rect 329 -279542 349 -275188
rect -350 -279570 349 -279542
rect -350 -279698 349 -279670
rect -350 -284052 265 -279698
rect 329 -284052 349 -279698
rect -350 -284080 349 -284052
rect -350 -284208 349 -284180
rect -350 -288562 265 -284208
rect 329 -288562 349 -284208
rect -350 -288590 349 -288562
<< via3 >>
rect 265 284208 329 288562
rect 265 279698 329 284052
rect 265 275188 329 279542
rect 265 270678 329 275032
rect 265 266168 329 270522
rect 265 261658 329 266012
rect 265 257148 329 261502
rect 265 252638 329 256992
rect 265 248128 329 252482
rect 265 243618 329 247972
rect 265 239108 329 243462
rect 265 234598 329 238952
rect 265 230088 329 234442
rect 265 225578 329 229932
rect 265 221068 329 225422
rect 265 216558 329 220912
rect 265 212048 329 216402
rect 265 207538 329 211892
rect 265 203028 329 207382
rect 265 198518 329 202872
rect 265 194008 329 198362
rect 265 189498 329 193852
rect 265 184988 329 189342
rect 265 180478 329 184832
rect 265 175968 329 180322
rect 265 171458 329 175812
rect 265 166948 329 171302
rect 265 162438 329 166792
rect 265 157928 329 162282
rect 265 153418 329 157772
rect 265 148908 329 153262
rect 265 144398 329 148752
rect 265 139888 329 144242
rect 265 135378 329 139732
rect 265 130868 329 135222
rect 265 126358 329 130712
rect 265 121848 329 126202
rect 265 117338 329 121692
rect 265 112828 329 117182
rect 265 108318 329 112672
rect 265 103808 329 108162
rect 265 99298 329 103652
rect 265 94788 329 99142
rect 265 90278 329 94632
rect 265 85768 329 90122
rect 265 81258 329 85612
rect 265 76748 329 81102
rect 265 72238 329 76592
rect 265 67728 329 72082
rect 265 63218 329 67572
rect 265 58708 329 63062
rect 265 54198 329 58552
rect 265 49688 329 54042
rect 265 45178 329 49532
rect 265 40668 329 45022
rect 265 36158 329 40512
rect 265 31648 329 36002
rect 265 27138 329 31492
rect 265 22628 329 26982
rect 265 18118 329 22472
rect 265 13608 329 17962
rect 265 9098 329 13452
rect 265 4588 329 8942
rect 265 78 329 4432
rect 265 -4432 329 -78
rect 265 -8942 329 -4588
rect 265 -13452 329 -9098
rect 265 -17962 329 -13608
rect 265 -22472 329 -18118
rect 265 -26982 329 -22628
rect 265 -31492 329 -27138
rect 265 -36002 329 -31648
rect 265 -40512 329 -36158
rect 265 -45022 329 -40668
rect 265 -49532 329 -45178
rect 265 -54042 329 -49688
rect 265 -58552 329 -54198
rect 265 -63062 329 -58708
rect 265 -67572 329 -63218
rect 265 -72082 329 -67728
rect 265 -76592 329 -72238
rect 265 -81102 329 -76748
rect 265 -85612 329 -81258
rect 265 -90122 329 -85768
rect 265 -94632 329 -90278
rect 265 -99142 329 -94788
rect 265 -103652 329 -99298
rect 265 -108162 329 -103808
rect 265 -112672 329 -108318
rect 265 -117182 329 -112828
rect 265 -121692 329 -117338
rect 265 -126202 329 -121848
rect 265 -130712 329 -126358
rect 265 -135222 329 -130868
rect 265 -139732 329 -135378
rect 265 -144242 329 -139888
rect 265 -148752 329 -144398
rect 265 -153262 329 -148908
rect 265 -157772 329 -153418
rect 265 -162282 329 -157928
rect 265 -166792 329 -162438
rect 265 -171302 329 -166948
rect 265 -175812 329 -171458
rect 265 -180322 329 -175968
rect 265 -184832 329 -180478
rect 265 -189342 329 -184988
rect 265 -193852 329 -189498
rect 265 -198362 329 -194008
rect 265 -202872 329 -198518
rect 265 -207382 329 -203028
rect 265 -211892 329 -207538
rect 265 -216402 329 -212048
rect 265 -220912 329 -216558
rect 265 -225422 329 -221068
rect 265 -229932 329 -225578
rect 265 -234442 329 -230088
rect 265 -238952 329 -234598
rect 265 -243462 329 -239108
rect 265 -247972 329 -243618
rect 265 -252482 329 -248128
rect 265 -256992 329 -252638
rect 265 -261502 329 -257148
rect 265 -266012 329 -261658
rect 265 -270522 329 -266168
rect 265 -275032 329 -270678
rect 265 -279542 329 -275188
rect 265 -284052 329 -279698
rect 265 -288562 329 -284208
<< mimcap >>
rect -250 288450 150 288490
rect -250 284320 -210 288450
rect 110 284320 150 288450
rect -250 284280 150 284320
rect -250 283940 150 283980
rect -250 279810 -210 283940
rect 110 279810 150 283940
rect -250 279770 150 279810
rect -250 279430 150 279470
rect -250 275300 -210 279430
rect 110 275300 150 279430
rect -250 275260 150 275300
rect -250 274920 150 274960
rect -250 270790 -210 274920
rect 110 270790 150 274920
rect -250 270750 150 270790
rect -250 270410 150 270450
rect -250 266280 -210 270410
rect 110 266280 150 270410
rect -250 266240 150 266280
rect -250 265900 150 265940
rect -250 261770 -210 265900
rect 110 261770 150 265900
rect -250 261730 150 261770
rect -250 261390 150 261430
rect -250 257260 -210 261390
rect 110 257260 150 261390
rect -250 257220 150 257260
rect -250 256880 150 256920
rect -250 252750 -210 256880
rect 110 252750 150 256880
rect -250 252710 150 252750
rect -250 252370 150 252410
rect -250 248240 -210 252370
rect 110 248240 150 252370
rect -250 248200 150 248240
rect -250 247860 150 247900
rect -250 243730 -210 247860
rect 110 243730 150 247860
rect -250 243690 150 243730
rect -250 243350 150 243390
rect -250 239220 -210 243350
rect 110 239220 150 243350
rect -250 239180 150 239220
rect -250 238840 150 238880
rect -250 234710 -210 238840
rect 110 234710 150 238840
rect -250 234670 150 234710
rect -250 234330 150 234370
rect -250 230200 -210 234330
rect 110 230200 150 234330
rect -250 230160 150 230200
rect -250 229820 150 229860
rect -250 225690 -210 229820
rect 110 225690 150 229820
rect -250 225650 150 225690
rect -250 225310 150 225350
rect -250 221180 -210 225310
rect 110 221180 150 225310
rect -250 221140 150 221180
rect -250 220800 150 220840
rect -250 216670 -210 220800
rect 110 216670 150 220800
rect -250 216630 150 216670
rect -250 216290 150 216330
rect -250 212160 -210 216290
rect 110 212160 150 216290
rect -250 212120 150 212160
rect -250 211780 150 211820
rect -250 207650 -210 211780
rect 110 207650 150 211780
rect -250 207610 150 207650
rect -250 207270 150 207310
rect -250 203140 -210 207270
rect 110 203140 150 207270
rect -250 203100 150 203140
rect -250 202760 150 202800
rect -250 198630 -210 202760
rect 110 198630 150 202760
rect -250 198590 150 198630
rect -250 198250 150 198290
rect -250 194120 -210 198250
rect 110 194120 150 198250
rect -250 194080 150 194120
rect -250 193740 150 193780
rect -250 189610 -210 193740
rect 110 189610 150 193740
rect -250 189570 150 189610
rect -250 189230 150 189270
rect -250 185100 -210 189230
rect 110 185100 150 189230
rect -250 185060 150 185100
rect -250 184720 150 184760
rect -250 180590 -210 184720
rect 110 180590 150 184720
rect -250 180550 150 180590
rect -250 180210 150 180250
rect -250 176080 -210 180210
rect 110 176080 150 180210
rect -250 176040 150 176080
rect -250 175700 150 175740
rect -250 171570 -210 175700
rect 110 171570 150 175700
rect -250 171530 150 171570
rect -250 171190 150 171230
rect -250 167060 -210 171190
rect 110 167060 150 171190
rect -250 167020 150 167060
rect -250 166680 150 166720
rect -250 162550 -210 166680
rect 110 162550 150 166680
rect -250 162510 150 162550
rect -250 162170 150 162210
rect -250 158040 -210 162170
rect 110 158040 150 162170
rect -250 158000 150 158040
rect -250 157660 150 157700
rect -250 153530 -210 157660
rect 110 153530 150 157660
rect -250 153490 150 153530
rect -250 153150 150 153190
rect -250 149020 -210 153150
rect 110 149020 150 153150
rect -250 148980 150 149020
rect -250 148640 150 148680
rect -250 144510 -210 148640
rect 110 144510 150 148640
rect -250 144470 150 144510
rect -250 144130 150 144170
rect -250 140000 -210 144130
rect 110 140000 150 144130
rect -250 139960 150 140000
rect -250 139620 150 139660
rect -250 135490 -210 139620
rect 110 135490 150 139620
rect -250 135450 150 135490
rect -250 135110 150 135150
rect -250 130980 -210 135110
rect 110 130980 150 135110
rect -250 130940 150 130980
rect -250 130600 150 130640
rect -250 126470 -210 130600
rect 110 126470 150 130600
rect -250 126430 150 126470
rect -250 126090 150 126130
rect -250 121960 -210 126090
rect 110 121960 150 126090
rect -250 121920 150 121960
rect -250 121580 150 121620
rect -250 117450 -210 121580
rect 110 117450 150 121580
rect -250 117410 150 117450
rect -250 117070 150 117110
rect -250 112940 -210 117070
rect 110 112940 150 117070
rect -250 112900 150 112940
rect -250 112560 150 112600
rect -250 108430 -210 112560
rect 110 108430 150 112560
rect -250 108390 150 108430
rect -250 108050 150 108090
rect -250 103920 -210 108050
rect 110 103920 150 108050
rect -250 103880 150 103920
rect -250 103540 150 103580
rect -250 99410 -210 103540
rect 110 99410 150 103540
rect -250 99370 150 99410
rect -250 99030 150 99070
rect -250 94900 -210 99030
rect 110 94900 150 99030
rect -250 94860 150 94900
rect -250 94520 150 94560
rect -250 90390 -210 94520
rect 110 90390 150 94520
rect -250 90350 150 90390
rect -250 90010 150 90050
rect -250 85880 -210 90010
rect 110 85880 150 90010
rect -250 85840 150 85880
rect -250 85500 150 85540
rect -250 81370 -210 85500
rect 110 81370 150 85500
rect -250 81330 150 81370
rect -250 80990 150 81030
rect -250 76860 -210 80990
rect 110 76860 150 80990
rect -250 76820 150 76860
rect -250 76480 150 76520
rect -250 72350 -210 76480
rect 110 72350 150 76480
rect -250 72310 150 72350
rect -250 71970 150 72010
rect -250 67840 -210 71970
rect 110 67840 150 71970
rect -250 67800 150 67840
rect -250 67460 150 67500
rect -250 63330 -210 67460
rect 110 63330 150 67460
rect -250 63290 150 63330
rect -250 62950 150 62990
rect -250 58820 -210 62950
rect 110 58820 150 62950
rect -250 58780 150 58820
rect -250 58440 150 58480
rect -250 54310 -210 58440
rect 110 54310 150 58440
rect -250 54270 150 54310
rect -250 53930 150 53970
rect -250 49800 -210 53930
rect 110 49800 150 53930
rect -250 49760 150 49800
rect -250 49420 150 49460
rect -250 45290 -210 49420
rect 110 45290 150 49420
rect -250 45250 150 45290
rect -250 44910 150 44950
rect -250 40780 -210 44910
rect 110 40780 150 44910
rect -250 40740 150 40780
rect -250 40400 150 40440
rect -250 36270 -210 40400
rect 110 36270 150 40400
rect -250 36230 150 36270
rect -250 35890 150 35930
rect -250 31760 -210 35890
rect 110 31760 150 35890
rect -250 31720 150 31760
rect -250 31380 150 31420
rect -250 27250 -210 31380
rect 110 27250 150 31380
rect -250 27210 150 27250
rect -250 26870 150 26910
rect -250 22740 -210 26870
rect 110 22740 150 26870
rect -250 22700 150 22740
rect -250 22360 150 22400
rect -250 18230 -210 22360
rect 110 18230 150 22360
rect -250 18190 150 18230
rect -250 17850 150 17890
rect -250 13720 -210 17850
rect 110 13720 150 17850
rect -250 13680 150 13720
rect -250 13340 150 13380
rect -250 9210 -210 13340
rect 110 9210 150 13340
rect -250 9170 150 9210
rect -250 8830 150 8870
rect -250 4700 -210 8830
rect 110 4700 150 8830
rect -250 4660 150 4700
rect -250 4320 150 4360
rect -250 190 -210 4320
rect 110 190 150 4320
rect -250 150 150 190
rect -250 -190 150 -150
rect -250 -4320 -210 -190
rect 110 -4320 150 -190
rect -250 -4360 150 -4320
rect -250 -4700 150 -4660
rect -250 -8830 -210 -4700
rect 110 -8830 150 -4700
rect -250 -8870 150 -8830
rect -250 -9210 150 -9170
rect -250 -13340 -210 -9210
rect 110 -13340 150 -9210
rect -250 -13380 150 -13340
rect -250 -13720 150 -13680
rect -250 -17850 -210 -13720
rect 110 -17850 150 -13720
rect -250 -17890 150 -17850
rect -250 -18230 150 -18190
rect -250 -22360 -210 -18230
rect 110 -22360 150 -18230
rect -250 -22400 150 -22360
rect -250 -22740 150 -22700
rect -250 -26870 -210 -22740
rect 110 -26870 150 -22740
rect -250 -26910 150 -26870
rect -250 -27250 150 -27210
rect -250 -31380 -210 -27250
rect 110 -31380 150 -27250
rect -250 -31420 150 -31380
rect -250 -31760 150 -31720
rect -250 -35890 -210 -31760
rect 110 -35890 150 -31760
rect -250 -35930 150 -35890
rect -250 -36270 150 -36230
rect -250 -40400 -210 -36270
rect 110 -40400 150 -36270
rect -250 -40440 150 -40400
rect -250 -40780 150 -40740
rect -250 -44910 -210 -40780
rect 110 -44910 150 -40780
rect -250 -44950 150 -44910
rect -250 -45290 150 -45250
rect -250 -49420 -210 -45290
rect 110 -49420 150 -45290
rect -250 -49460 150 -49420
rect -250 -49800 150 -49760
rect -250 -53930 -210 -49800
rect 110 -53930 150 -49800
rect -250 -53970 150 -53930
rect -250 -54310 150 -54270
rect -250 -58440 -210 -54310
rect 110 -58440 150 -54310
rect -250 -58480 150 -58440
rect -250 -58820 150 -58780
rect -250 -62950 -210 -58820
rect 110 -62950 150 -58820
rect -250 -62990 150 -62950
rect -250 -63330 150 -63290
rect -250 -67460 -210 -63330
rect 110 -67460 150 -63330
rect -250 -67500 150 -67460
rect -250 -67840 150 -67800
rect -250 -71970 -210 -67840
rect 110 -71970 150 -67840
rect -250 -72010 150 -71970
rect -250 -72350 150 -72310
rect -250 -76480 -210 -72350
rect 110 -76480 150 -72350
rect -250 -76520 150 -76480
rect -250 -76860 150 -76820
rect -250 -80990 -210 -76860
rect 110 -80990 150 -76860
rect -250 -81030 150 -80990
rect -250 -81370 150 -81330
rect -250 -85500 -210 -81370
rect 110 -85500 150 -81370
rect -250 -85540 150 -85500
rect -250 -85880 150 -85840
rect -250 -90010 -210 -85880
rect 110 -90010 150 -85880
rect -250 -90050 150 -90010
rect -250 -90390 150 -90350
rect -250 -94520 -210 -90390
rect 110 -94520 150 -90390
rect -250 -94560 150 -94520
rect -250 -94900 150 -94860
rect -250 -99030 -210 -94900
rect 110 -99030 150 -94900
rect -250 -99070 150 -99030
rect -250 -99410 150 -99370
rect -250 -103540 -210 -99410
rect 110 -103540 150 -99410
rect -250 -103580 150 -103540
rect -250 -103920 150 -103880
rect -250 -108050 -210 -103920
rect 110 -108050 150 -103920
rect -250 -108090 150 -108050
rect -250 -108430 150 -108390
rect -250 -112560 -210 -108430
rect 110 -112560 150 -108430
rect -250 -112600 150 -112560
rect -250 -112940 150 -112900
rect -250 -117070 -210 -112940
rect 110 -117070 150 -112940
rect -250 -117110 150 -117070
rect -250 -117450 150 -117410
rect -250 -121580 -210 -117450
rect 110 -121580 150 -117450
rect -250 -121620 150 -121580
rect -250 -121960 150 -121920
rect -250 -126090 -210 -121960
rect 110 -126090 150 -121960
rect -250 -126130 150 -126090
rect -250 -126470 150 -126430
rect -250 -130600 -210 -126470
rect 110 -130600 150 -126470
rect -250 -130640 150 -130600
rect -250 -130980 150 -130940
rect -250 -135110 -210 -130980
rect 110 -135110 150 -130980
rect -250 -135150 150 -135110
rect -250 -135490 150 -135450
rect -250 -139620 -210 -135490
rect 110 -139620 150 -135490
rect -250 -139660 150 -139620
rect -250 -140000 150 -139960
rect -250 -144130 -210 -140000
rect 110 -144130 150 -140000
rect -250 -144170 150 -144130
rect -250 -144510 150 -144470
rect -250 -148640 -210 -144510
rect 110 -148640 150 -144510
rect -250 -148680 150 -148640
rect -250 -149020 150 -148980
rect -250 -153150 -210 -149020
rect 110 -153150 150 -149020
rect -250 -153190 150 -153150
rect -250 -153530 150 -153490
rect -250 -157660 -210 -153530
rect 110 -157660 150 -153530
rect -250 -157700 150 -157660
rect -250 -158040 150 -158000
rect -250 -162170 -210 -158040
rect 110 -162170 150 -158040
rect -250 -162210 150 -162170
rect -250 -162550 150 -162510
rect -250 -166680 -210 -162550
rect 110 -166680 150 -162550
rect -250 -166720 150 -166680
rect -250 -167060 150 -167020
rect -250 -171190 -210 -167060
rect 110 -171190 150 -167060
rect -250 -171230 150 -171190
rect -250 -171570 150 -171530
rect -250 -175700 -210 -171570
rect 110 -175700 150 -171570
rect -250 -175740 150 -175700
rect -250 -176080 150 -176040
rect -250 -180210 -210 -176080
rect 110 -180210 150 -176080
rect -250 -180250 150 -180210
rect -250 -180590 150 -180550
rect -250 -184720 -210 -180590
rect 110 -184720 150 -180590
rect -250 -184760 150 -184720
rect -250 -185100 150 -185060
rect -250 -189230 -210 -185100
rect 110 -189230 150 -185100
rect -250 -189270 150 -189230
rect -250 -189610 150 -189570
rect -250 -193740 -210 -189610
rect 110 -193740 150 -189610
rect -250 -193780 150 -193740
rect -250 -194120 150 -194080
rect -250 -198250 -210 -194120
rect 110 -198250 150 -194120
rect -250 -198290 150 -198250
rect -250 -198630 150 -198590
rect -250 -202760 -210 -198630
rect 110 -202760 150 -198630
rect -250 -202800 150 -202760
rect -250 -203140 150 -203100
rect -250 -207270 -210 -203140
rect 110 -207270 150 -203140
rect -250 -207310 150 -207270
rect -250 -207650 150 -207610
rect -250 -211780 -210 -207650
rect 110 -211780 150 -207650
rect -250 -211820 150 -211780
rect -250 -212160 150 -212120
rect -250 -216290 -210 -212160
rect 110 -216290 150 -212160
rect -250 -216330 150 -216290
rect -250 -216670 150 -216630
rect -250 -220800 -210 -216670
rect 110 -220800 150 -216670
rect -250 -220840 150 -220800
rect -250 -221180 150 -221140
rect -250 -225310 -210 -221180
rect 110 -225310 150 -221180
rect -250 -225350 150 -225310
rect -250 -225690 150 -225650
rect -250 -229820 -210 -225690
rect 110 -229820 150 -225690
rect -250 -229860 150 -229820
rect -250 -230200 150 -230160
rect -250 -234330 -210 -230200
rect 110 -234330 150 -230200
rect -250 -234370 150 -234330
rect -250 -234710 150 -234670
rect -250 -238840 -210 -234710
rect 110 -238840 150 -234710
rect -250 -238880 150 -238840
rect -250 -239220 150 -239180
rect -250 -243350 -210 -239220
rect 110 -243350 150 -239220
rect -250 -243390 150 -243350
rect -250 -243730 150 -243690
rect -250 -247860 -210 -243730
rect 110 -247860 150 -243730
rect -250 -247900 150 -247860
rect -250 -248240 150 -248200
rect -250 -252370 -210 -248240
rect 110 -252370 150 -248240
rect -250 -252410 150 -252370
rect -250 -252750 150 -252710
rect -250 -256880 -210 -252750
rect 110 -256880 150 -252750
rect -250 -256920 150 -256880
rect -250 -257260 150 -257220
rect -250 -261390 -210 -257260
rect 110 -261390 150 -257260
rect -250 -261430 150 -261390
rect -250 -261770 150 -261730
rect -250 -265900 -210 -261770
rect 110 -265900 150 -261770
rect -250 -265940 150 -265900
rect -250 -266280 150 -266240
rect -250 -270410 -210 -266280
rect 110 -270410 150 -266280
rect -250 -270450 150 -270410
rect -250 -270790 150 -270750
rect -250 -274920 -210 -270790
rect 110 -274920 150 -270790
rect -250 -274960 150 -274920
rect -250 -275300 150 -275260
rect -250 -279430 -210 -275300
rect 110 -279430 150 -275300
rect -250 -279470 150 -279430
rect -250 -279810 150 -279770
rect -250 -283940 -210 -279810
rect 110 -283940 150 -279810
rect -250 -283980 150 -283940
rect -250 -284320 150 -284280
rect -250 -288450 -210 -284320
rect 110 -288450 150 -284320
rect -250 -288490 150 -288450
<< mimcapcontact >>
rect -210 284320 110 288450
rect -210 279810 110 283940
rect -210 275300 110 279430
rect -210 270790 110 274920
rect -210 266280 110 270410
rect -210 261770 110 265900
rect -210 257260 110 261390
rect -210 252750 110 256880
rect -210 248240 110 252370
rect -210 243730 110 247860
rect -210 239220 110 243350
rect -210 234710 110 238840
rect -210 230200 110 234330
rect -210 225690 110 229820
rect -210 221180 110 225310
rect -210 216670 110 220800
rect -210 212160 110 216290
rect -210 207650 110 211780
rect -210 203140 110 207270
rect -210 198630 110 202760
rect -210 194120 110 198250
rect -210 189610 110 193740
rect -210 185100 110 189230
rect -210 180590 110 184720
rect -210 176080 110 180210
rect -210 171570 110 175700
rect -210 167060 110 171190
rect -210 162550 110 166680
rect -210 158040 110 162170
rect -210 153530 110 157660
rect -210 149020 110 153150
rect -210 144510 110 148640
rect -210 140000 110 144130
rect -210 135490 110 139620
rect -210 130980 110 135110
rect -210 126470 110 130600
rect -210 121960 110 126090
rect -210 117450 110 121580
rect -210 112940 110 117070
rect -210 108430 110 112560
rect -210 103920 110 108050
rect -210 99410 110 103540
rect -210 94900 110 99030
rect -210 90390 110 94520
rect -210 85880 110 90010
rect -210 81370 110 85500
rect -210 76860 110 80990
rect -210 72350 110 76480
rect -210 67840 110 71970
rect -210 63330 110 67460
rect -210 58820 110 62950
rect -210 54310 110 58440
rect -210 49800 110 53930
rect -210 45290 110 49420
rect -210 40780 110 44910
rect -210 36270 110 40400
rect -210 31760 110 35890
rect -210 27250 110 31380
rect -210 22740 110 26870
rect -210 18230 110 22360
rect -210 13720 110 17850
rect -210 9210 110 13340
rect -210 4700 110 8830
rect -210 190 110 4320
rect -210 -4320 110 -190
rect -210 -8830 110 -4700
rect -210 -13340 110 -9210
rect -210 -17850 110 -13720
rect -210 -22360 110 -18230
rect -210 -26870 110 -22740
rect -210 -31380 110 -27250
rect -210 -35890 110 -31760
rect -210 -40400 110 -36270
rect -210 -44910 110 -40780
rect -210 -49420 110 -45290
rect -210 -53930 110 -49800
rect -210 -58440 110 -54310
rect -210 -62950 110 -58820
rect -210 -67460 110 -63330
rect -210 -71970 110 -67840
rect -210 -76480 110 -72350
rect -210 -80990 110 -76860
rect -210 -85500 110 -81370
rect -210 -90010 110 -85880
rect -210 -94520 110 -90390
rect -210 -99030 110 -94900
rect -210 -103540 110 -99410
rect -210 -108050 110 -103920
rect -210 -112560 110 -108430
rect -210 -117070 110 -112940
rect -210 -121580 110 -117450
rect -210 -126090 110 -121960
rect -210 -130600 110 -126470
rect -210 -135110 110 -130980
rect -210 -139620 110 -135490
rect -210 -144130 110 -140000
rect -210 -148640 110 -144510
rect -210 -153150 110 -149020
rect -210 -157660 110 -153530
rect -210 -162170 110 -158040
rect -210 -166680 110 -162550
rect -210 -171190 110 -167060
rect -210 -175700 110 -171570
rect -210 -180210 110 -176080
rect -210 -184720 110 -180590
rect -210 -189230 110 -185100
rect -210 -193740 110 -189610
rect -210 -198250 110 -194120
rect -210 -202760 110 -198630
rect -210 -207270 110 -203140
rect -210 -211780 110 -207650
rect -210 -216290 110 -212160
rect -210 -220800 110 -216670
rect -210 -225310 110 -221180
rect -210 -229820 110 -225690
rect -210 -234330 110 -230200
rect -210 -238840 110 -234710
rect -210 -243350 110 -239220
rect -210 -247860 110 -243730
rect -210 -252370 110 -248240
rect -210 -256880 110 -252750
rect -210 -261390 110 -257260
rect -210 -265900 110 -261770
rect -210 -270410 110 -266280
rect -210 -274920 110 -270790
rect -210 -279430 110 -275300
rect -210 -283940 110 -279810
rect -210 -288450 110 -284320
<< metal4 >>
rect -102 288451 2 288640
rect 218 288578 322 288640
rect 218 288562 345 288578
rect -211 288450 111 288451
rect -211 284320 -210 288450
rect 110 284320 111 288450
rect -211 284319 111 284320
rect -102 283941 2 284319
rect 218 284208 265 288562
rect 329 284208 345 288562
rect 218 284192 345 284208
rect 218 284068 322 284192
rect 218 284052 345 284068
rect -211 283940 111 283941
rect -211 279810 -210 283940
rect 110 279810 111 283940
rect -211 279809 111 279810
rect -102 279431 2 279809
rect 218 279698 265 284052
rect 329 279698 345 284052
rect 218 279682 345 279698
rect 218 279558 322 279682
rect 218 279542 345 279558
rect -211 279430 111 279431
rect -211 275300 -210 279430
rect 110 275300 111 279430
rect -211 275299 111 275300
rect -102 274921 2 275299
rect 218 275188 265 279542
rect 329 275188 345 279542
rect 218 275172 345 275188
rect 218 275048 322 275172
rect 218 275032 345 275048
rect -211 274920 111 274921
rect -211 270790 -210 274920
rect 110 270790 111 274920
rect -211 270789 111 270790
rect -102 270411 2 270789
rect 218 270678 265 275032
rect 329 270678 345 275032
rect 218 270662 345 270678
rect 218 270538 322 270662
rect 218 270522 345 270538
rect -211 270410 111 270411
rect -211 266280 -210 270410
rect 110 266280 111 270410
rect -211 266279 111 266280
rect -102 265901 2 266279
rect 218 266168 265 270522
rect 329 266168 345 270522
rect 218 266152 345 266168
rect 218 266028 322 266152
rect 218 266012 345 266028
rect -211 265900 111 265901
rect -211 261770 -210 265900
rect 110 261770 111 265900
rect -211 261769 111 261770
rect -102 261391 2 261769
rect 218 261658 265 266012
rect 329 261658 345 266012
rect 218 261642 345 261658
rect 218 261518 322 261642
rect 218 261502 345 261518
rect -211 261390 111 261391
rect -211 257260 -210 261390
rect 110 257260 111 261390
rect -211 257259 111 257260
rect -102 256881 2 257259
rect 218 257148 265 261502
rect 329 257148 345 261502
rect 218 257132 345 257148
rect 218 257008 322 257132
rect 218 256992 345 257008
rect -211 256880 111 256881
rect -211 252750 -210 256880
rect 110 252750 111 256880
rect -211 252749 111 252750
rect -102 252371 2 252749
rect 218 252638 265 256992
rect 329 252638 345 256992
rect 218 252622 345 252638
rect 218 252498 322 252622
rect 218 252482 345 252498
rect -211 252370 111 252371
rect -211 248240 -210 252370
rect 110 248240 111 252370
rect -211 248239 111 248240
rect -102 247861 2 248239
rect 218 248128 265 252482
rect 329 248128 345 252482
rect 218 248112 345 248128
rect 218 247988 322 248112
rect 218 247972 345 247988
rect -211 247860 111 247861
rect -211 243730 -210 247860
rect 110 243730 111 247860
rect -211 243729 111 243730
rect -102 243351 2 243729
rect 218 243618 265 247972
rect 329 243618 345 247972
rect 218 243602 345 243618
rect 218 243478 322 243602
rect 218 243462 345 243478
rect -211 243350 111 243351
rect -211 239220 -210 243350
rect 110 239220 111 243350
rect -211 239219 111 239220
rect -102 238841 2 239219
rect 218 239108 265 243462
rect 329 239108 345 243462
rect 218 239092 345 239108
rect 218 238968 322 239092
rect 218 238952 345 238968
rect -211 238840 111 238841
rect -211 234710 -210 238840
rect 110 234710 111 238840
rect -211 234709 111 234710
rect -102 234331 2 234709
rect 218 234598 265 238952
rect 329 234598 345 238952
rect 218 234582 345 234598
rect 218 234458 322 234582
rect 218 234442 345 234458
rect -211 234330 111 234331
rect -211 230200 -210 234330
rect 110 230200 111 234330
rect -211 230199 111 230200
rect -102 229821 2 230199
rect 218 230088 265 234442
rect 329 230088 345 234442
rect 218 230072 345 230088
rect 218 229948 322 230072
rect 218 229932 345 229948
rect -211 229820 111 229821
rect -211 225690 -210 229820
rect 110 225690 111 229820
rect -211 225689 111 225690
rect -102 225311 2 225689
rect 218 225578 265 229932
rect 329 225578 345 229932
rect 218 225562 345 225578
rect 218 225438 322 225562
rect 218 225422 345 225438
rect -211 225310 111 225311
rect -211 221180 -210 225310
rect 110 221180 111 225310
rect -211 221179 111 221180
rect -102 220801 2 221179
rect 218 221068 265 225422
rect 329 221068 345 225422
rect 218 221052 345 221068
rect 218 220928 322 221052
rect 218 220912 345 220928
rect -211 220800 111 220801
rect -211 216670 -210 220800
rect 110 216670 111 220800
rect -211 216669 111 216670
rect -102 216291 2 216669
rect 218 216558 265 220912
rect 329 216558 345 220912
rect 218 216542 345 216558
rect 218 216418 322 216542
rect 218 216402 345 216418
rect -211 216290 111 216291
rect -211 212160 -210 216290
rect 110 212160 111 216290
rect -211 212159 111 212160
rect -102 211781 2 212159
rect 218 212048 265 216402
rect 329 212048 345 216402
rect 218 212032 345 212048
rect 218 211908 322 212032
rect 218 211892 345 211908
rect -211 211780 111 211781
rect -211 207650 -210 211780
rect 110 207650 111 211780
rect -211 207649 111 207650
rect -102 207271 2 207649
rect 218 207538 265 211892
rect 329 207538 345 211892
rect 218 207522 345 207538
rect 218 207398 322 207522
rect 218 207382 345 207398
rect -211 207270 111 207271
rect -211 203140 -210 207270
rect 110 203140 111 207270
rect -211 203139 111 203140
rect -102 202761 2 203139
rect 218 203028 265 207382
rect 329 203028 345 207382
rect 218 203012 345 203028
rect 218 202888 322 203012
rect 218 202872 345 202888
rect -211 202760 111 202761
rect -211 198630 -210 202760
rect 110 198630 111 202760
rect -211 198629 111 198630
rect -102 198251 2 198629
rect 218 198518 265 202872
rect 329 198518 345 202872
rect 218 198502 345 198518
rect 218 198378 322 198502
rect 218 198362 345 198378
rect -211 198250 111 198251
rect -211 194120 -210 198250
rect 110 194120 111 198250
rect -211 194119 111 194120
rect -102 193741 2 194119
rect 218 194008 265 198362
rect 329 194008 345 198362
rect 218 193992 345 194008
rect 218 193868 322 193992
rect 218 193852 345 193868
rect -211 193740 111 193741
rect -211 189610 -210 193740
rect 110 189610 111 193740
rect -211 189609 111 189610
rect -102 189231 2 189609
rect 218 189498 265 193852
rect 329 189498 345 193852
rect 218 189482 345 189498
rect 218 189358 322 189482
rect 218 189342 345 189358
rect -211 189230 111 189231
rect -211 185100 -210 189230
rect 110 185100 111 189230
rect -211 185099 111 185100
rect -102 184721 2 185099
rect 218 184988 265 189342
rect 329 184988 345 189342
rect 218 184972 345 184988
rect 218 184848 322 184972
rect 218 184832 345 184848
rect -211 184720 111 184721
rect -211 180590 -210 184720
rect 110 180590 111 184720
rect -211 180589 111 180590
rect -102 180211 2 180589
rect 218 180478 265 184832
rect 329 180478 345 184832
rect 218 180462 345 180478
rect 218 180338 322 180462
rect 218 180322 345 180338
rect -211 180210 111 180211
rect -211 176080 -210 180210
rect 110 176080 111 180210
rect -211 176079 111 176080
rect -102 175701 2 176079
rect 218 175968 265 180322
rect 329 175968 345 180322
rect 218 175952 345 175968
rect 218 175828 322 175952
rect 218 175812 345 175828
rect -211 175700 111 175701
rect -211 171570 -210 175700
rect 110 171570 111 175700
rect -211 171569 111 171570
rect -102 171191 2 171569
rect 218 171458 265 175812
rect 329 171458 345 175812
rect 218 171442 345 171458
rect 218 171318 322 171442
rect 218 171302 345 171318
rect -211 171190 111 171191
rect -211 167060 -210 171190
rect 110 167060 111 171190
rect -211 167059 111 167060
rect -102 166681 2 167059
rect 218 166948 265 171302
rect 329 166948 345 171302
rect 218 166932 345 166948
rect 218 166808 322 166932
rect 218 166792 345 166808
rect -211 166680 111 166681
rect -211 162550 -210 166680
rect 110 162550 111 166680
rect -211 162549 111 162550
rect -102 162171 2 162549
rect 218 162438 265 166792
rect 329 162438 345 166792
rect 218 162422 345 162438
rect 218 162298 322 162422
rect 218 162282 345 162298
rect -211 162170 111 162171
rect -211 158040 -210 162170
rect 110 158040 111 162170
rect -211 158039 111 158040
rect -102 157661 2 158039
rect 218 157928 265 162282
rect 329 157928 345 162282
rect 218 157912 345 157928
rect 218 157788 322 157912
rect 218 157772 345 157788
rect -211 157660 111 157661
rect -211 153530 -210 157660
rect 110 153530 111 157660
rect -211 153529 111 153530
rect -102 153151 2 153529
rect 218 153418 265 157772
rect 329 153418 345 157772
rect 218 153402 345 153418
rect 218 153278 322 153402
rect 218 153262 345 153278
rect -211 153150 111 153151
rect -211 149020 -210 153150
rect 110 149020 111 153150
rect -211 149019 111 149020
rect -102 148641 2 149019
rect 218 148908 265 153262
rect 329 148908 345 153262
rect 218 148892 345 148908
rect 218 148768 322 148892
rect 218 148752 345 148768
rect -211 148640 111 148641
rect -211 144510 -210 148640
rect 110 144510 111 148640
rect -211 144509 111 144510
rect -102 144131 2 144509
rect 218 144398 265 148752
rect 329 144398 345 148752
rect 218 144382 345 144398
rect 218 144258 322 144382
rect 218 144242 345 144258
rect -211 144130 111 144131
rect -211 140000 -210 144130
rect 110 140000 111 144130
rect -211 139999 111 140000
rect -102 139621 2 139999
rect 218 139888 265 144242
rect 329 139888 345 144242
rect 218 139872 345 139888
rect 218 139748 322 139872
rect 218 139732 345 139748
rect -211 139620 111 139621
rect -211 135490 -210 139620
rect 110 135490 111 139620
rect -211 135489 111 135490
rect -102 135111 2 135489
rect 218 135378 265 139732
rect 329 135378 345 139732
rect 218 135362 345 135378
rect 218 135238 322 135362
rect 218 135222 345 135238
rect -211 135110 111 135111
rect -211 130980 -210 135110
rect 110 130980 111 135110
rect -211 130979 111 130980
rect -102 130601 2 130979
rect 218 130868 265 135222
rect 329 130868 345 135222
rect 218 130852 345 130868
rect 218 130728 322 130852
rect 218 130712 345 130728
rect -211 130600 111 130601
rect -211 126470 -210 130600
rect 110 126470 111 130600
rect -211 126469 111 126470
rect -102 126091 2 126469
rect 218 126358 265 130712
rect 329 126358 345 130712
rect 218 126342 345 126358
rect 218 126218 322 126342
rect 218 126202 345 126218
rect -211 126090 111 126091
rect -211 121960 -210 126090
rect 110 121960 111 126090
rect -211 121959 111 121960
rect -102 121581 2 121959
rect 218 121848 265 126202
rect 329 121848 345 126202
rect 218 121832 345 121848
rect 218 121708 322 121832
rect 218 121692 345 121708
rect -211 121580 111 121581
rect -211 117450 -210 121580
rect 110 117450 111 121580
rect -211 117449 111 117450
rect -102 117071 2 117449
rect 218 117338 265 121692
rect 329 117338 345 121692
rect 218 117322 345 117338
rect 218 117198 322 117322
rect 218 117182 345 117198
rect -211 117070 111 117071
rect -211 112940 -210 117070
rect 110 112940 111 117070
rect -211 112939 111 112940
rect -102 112561 2 112939
rect 218 112828 265 117182
rect 329 112828 345 117182
rect 218 112812 345 112828
rect 218 112688 322 112812
rect 218 112672 345 112688
rect -211 112560 111 112561
rect -211 108430 -210 112560
rect 110 108430 111 112560
rect -211 108429 111 108430
rect -102 108051 2 108429
rect 218 108318 265 112672
rect 329 108318 345 112672
rect 218 108302 345 108318
rect 218 108178 322 108302
rect 218 108162 345 108178
rect -211 108050 111 108051
rect -211 103920 -210 108050
rect 110 103920 111 108050
rect -211 103919 111 103920
rect -102 103541 2 103919
rect 218 103808 265 108162
rect 329 103808 345 108162
rect 218 103792 345 103808
rect 218 103668 322 103792
rect 218 103652 345 103668
rect -211 103540 111 103541
rect -211 99410 -210 103540
rect 110 99410 111 103540
rect -211 99409 111 99410
rect -102 99031 2 99409
rect 218 99298 265 103652
rect 329 99298 345 103652
rect 218 99282 345 99298
rect 218 99158 322 99282
rect 218 99142 345 99158
rect -211 99030 111 99031
rect -211 94900 -210 99030
rect 110 94900 111 99030
rect -211 94899 111 94900
rect -102 94521 2 94899
rect 218 94788 265 99142
rect 329 94788 345 99142
rect 218 94772 345 94788
rect 218 94648 322 94772
rect 218 94632 345 94648
rect -211 94520 111 94521
rect -211 90390 -210 94520
rect 110 90390 111 94520
rect -211 90389 111 90390
rect -102 90011 2 90389
rect 218 90278 265 94632
rect 329 90278 345 94632
rect 218 90262 345 90278
rect 218 90138 322 90262
rect 218 90122 345 90138
rect -211 90010 111 90011
rect -211 85880 -210 90010
rect 110 85880 111 90010
rect -211 85879 111 85880
rect -102 85501 2 85879
rect 218 85768 265 90122
rect 329 85768 345 90122
rect 218 85752 345 85768
rect 218 85628 322 85752
rect 218 85612 345 85628
rect -211 85500 111 85501
rect -211 81370 -210 85500
rect 110 81370 111 85500
rect -211 81369 111 81370
rect -102 80991 2 81369
rect 218 81258 265 85612
rect 329 81258 345 85612
rect 218 81242 345 81258
rect 218 81118 322 81242
rect 218 81102 345 81118
rect -211 80990 111 80991
rect -211 76860 -210 80990
rect 110 76860 111 80990
rect -211 76859 111 76860
rect -102 76481 2 76859
rect 218 76748 265 81102
rect 329 76748 345 81102
rect 218 76732 345 76748
rect 218 76608 322 76732
rect 218 76592 345 76608
rect -211 76480 111 76481
rect -211 72350 -210 76480
rect 110 72350 111 76480
rect -211 72349 111 72350
rect -102 71971 2 72349
rect 218 72238 265 76592
rect 329 72238 345 76592
rect 218 72222 345 72238
rect 218 72098 322 72222
rect 218 72082 345 72098
rect -211 71970 111 71971
rect -211 67840 -210 71970
rect 110 67840 111 71970
rect -211 67839 111 67840
rect -102 67461 2 67839
rect 218 67728 265 72082
rect 329 67728 345 72082
rect 218 67712 345 67728
rect 218 67588 322 67712
rect 218 67572 345 67588
rect -211 67460 111 67461
rect -211 63330 -210 67460
rect 110 63330 111 67460
rect -211 63329 111 63330
rect -102 62951 2 63329
rect 218 63218 265 67572
rect 329 63218 345 67572
rect 218 63202 345 63218
rect 218 63078 322 63202
rect 218 63062 345 63078
rect -211 62950 111 62951
rect -211 58820 -210 62950
rect 110 58820 111 62950
rect -211 58819 111 58820
rect -102 58441 2 58819
rect 218 58708 265 63062
rect 329 58708 345 63062
rect 218 58692 345 58708
rect 218 58568 322 58692
rect 218 58552 345 58568
rect -211 58440 111 58441
rect -211 54310 -210 58440
rect 110 54310 111 58440
rect -211 54309 111 54310
rect -102 53931 2 54309
rect 218 54198 265 58552
rect 329 54198 345 58552
rect 218 54182 345 54198
rect 218 54058 322 54182
rect 218 54042 345 54058
rect -211 53930 111 53931
rect -211 49800 -210 53930
rect 110 49800 111 53930
rect -211 49799 111 49800
rect -102 49421 2 49799
rect 218 49688 265 54042
rect 329 49688 345 54042
rect 218 49672 345 49688
rect 218 49548 322 49672
rect 218 49532 345 49548
rect -211 49420 111 49421
rect -211 45290 -210 49420
rect 110 45290 111 49420
rect -211 45289 111 45290
rect -102 44911 2 45289
rect 218 45178 265 49532
rect 329 45178 345 49532
rect 218 45162 345 45178
rect 218 45038 322 45162
rect 218 45022 345 45038
rect -211 44910 111 44911
rect -211 40780 -210 44910
rect 110 40780 111 44910
rect -211 40779 111 40780
rect -102 40401 2 40779
rect 218 40668 265 45022
rect 329 40668 345 45022
rect 218 40652 345 40668
rect 218 40528 322 40652
rect 218 40512 345 40528
rect -211 40400 111 40401
rect -211 36270 -210 40400
rect 110 36270 111 40400
rect -211 36269 111 36270
rect -102 35891 2 36269
rect 218 36158 265 40512
rect 329 36158 345 40512
rect 218 36142 345 36158
rect 218 36018 322 36142
rect 218 36002 345 36018
rect -211 35890 111 35891
rect -211 31760 -210 35890
rect 110 31760 111 35890
rect -211 31759 111 31760
rect -102 31381 2 31759
rect 218 31648 265 36002
rect 329 31648 345 36002
rect 218 31632 345 31648
rect 218 31508 322 31632
rect 218 31492 345 31508
rect -211 31380 111 31381
rect -211 27250 -210 31380
rect 110 27250 111 31380
rect -211 27249 111 27250
rect -102 26871 2 27249
rect 218 27138 265 31492
rect 329 27138 345 31492
rect 218 27122 345 27138
rect 218 26998 322 27122
rect 218 26982 345 26998
rect -211 26870 111 26871
rect -211 22740 -210 26870
rect 110 22740 111 26870
rect -211 22739 111 22740
rect -102 22361 2 22739
rect 218 22628 265 26982
rect 329 22628 345 26982
rect 218 22612 345 22628
rect 218 22488 322 22612
rect 218 22472 345 22488
rect -211 22360 111 22361
rect -211 18230 -210 22360
rect 110 18230 111 22360
rect -211 18229 111 18230
rect -102 17851 2 18229
rect 218 18118 265 22472
rect 329 18118 345 22472
rect 218 18102 345 18118
rect 218 17978 322 18102
rect 218 17962 345 17978
rect -211 17850 111 17851
rect -211 13720 -210 17850
rect 110 13720 111 17850
rect -211 13719 111 13720
rect -102 13341 2 13719
rect 218 13608 265 17962
rect 329 13608 345 17962
rect 218 13592 345 13608
rect 218 13468 322 13592
rect 218 13452 345 13468
rect -211 13340 111 13341
rect -211 9210 -210 13340
rect 110 9210 111 13340
rect -211 9209 111 9210
rect -102 8831 2 9209
rect 218 9098 265 13452
rect 329 9098 345 13452
rect 218 9082 345 9098
rect 218 8958 322 9082
rect 218 8942 345 8958
rect -211 8830 111 8831
rect -211 4700 -210 8830
rect 110 4700 111 8830
rect -211 4699 111 4700
rect -102 4321 2 4699
rect 218 4588 265 8942
rect 329 4588 345 8942
rect 218 4572 345 4588
rect 218 4448 322 4572
rect 218 4432 345 4448
rect -211 4320 111 4321
rect -211 190 -210 4320
rect 110 190 111 4320
rect -211 189 111 190
rect -102 -189 2 189
rect 218 78 265 4432
rect 329 78 345 4432
rect 218 62 345 78
rect 218 -62 322 62
rect 218 -78 345 -62
rect -211 -190 111 -189
rect -211 -4320 -210 -190
rect 110 -4320 111 -190
rect -211 -4321 111 -4320
rect -102 -4699 2 -4321
rect 218 -4432 265 -78
rect 329 -4432 345 -78
rect 218 -4448 345 -4432
rect 218 -4572 322 -4448
rect 218 -4588 345 -4572
rect -211 -4700 111 -4699
rect -211 -8830 -210 -4700
rect 110 -8830 111 -4700
rect -211 -8831 111 -8830
rect -102 -9209 2 -8831
rect 218 -8942 265 -4588
rect 329 -8942 345 -4588
rect 218 -8958 345 -8942
rect 218 -9082 322 -8958
rect 218 -9098 345 -9082
rect -211 -9210 111 -9209
rect -211 -13340 -210 -9210
rect 110 -13340 111 -9210
rect -211 -13341 111 -13340
rect -102 -13719 2 -13341
rect 218 -13452 265 -9098
rect 329 -13452 345 -9098
rect 218 -13468 345 -13452
rect 218 -13592 322 -13468
rect 218 -13608 345 -13592
rect -211 -13720 111 -13719
rect -211 -17850 -210 -13720
rect 110 -17850 111 -13720
rect -211 -17851 111 -17850
rect -102 -18229 2 -17851
rect 218 -17962 265 -13608
rect 329 -17962 345 -13608
rect 218 -17978 345 -17962
rect 218 -18102 322 -17978
rect 218 -18118 345 -18102
rect -211 -18230 111 -18229
rect -211 -22360 -210 -18230
rect 110 -22360 111 -18230
rect -211 -22361 111 -22360
rect -102 -22739 2 -22361
rect 218 -22472 265 -18118
rect 329 -22472 345 -18118
rect 218 -22488 345 -22472
rect 218 -22612 322 -22488
rect 218 -22628 345 -22612
rect -211 -22740 111 -22739
rect -211 -26870 -210 -22740
rect 110 -26870 111 -22740
rect -211 -26871 111 -26870
rect -102 -27249 2 -26871
rect 218 -26982 265 -22628
rect 329 -26982 345 -22628
rect 218 -26998 345 -26982
rect 218 -27122 322 -26998
rect 218 -27138 345 -27122
rect -211 -27250 111 -27249
rect -211 -31380 -210 -27250
rect 110 -31380 111 -27250
rect -211 -31381 111 -31380
rect -102 -31759 2 -31381
rect 218 -31492 265 -27138
rect 329 -31492 345 -27138
rect 218 -31508 345 -31492
rect 218 -31632 322 -31508
rect 218 -31648 345 -31632
rect -211 -31760 111 -31759
rect -211 -35890 -210 -31760
rect 110 -35890 111 -31760
rect -211 -35891 111 -35890
rect -102 -36269 2 -35891
rect 218 -36002 265 -31648
rect 329 -36002 345 -31648
rect 218 -36018 345 -36002
rect 218 -36142 322 -36018
rect 218 -36158 345 -36142
rect -211 -36270 111 -36269
rect -211 -40400 -210 -36270
rect 110 -40400 111 -36270
rect -211 -40401 111 -40400
rect -102 -40779 2 -40401
rect 218 -40512 265 -36158
rect 329 -40512 345 -36158
rect 218 -40528 345 -40512
rect 218 -40652 322 -40528
rect 218 -40668 345 -40652
rect -211 -40780 111 -40779
rect -211 -44910 -210 -40780
rect 110 -44910 111 -40780
rect -211 -44911 111 -44910
rect -102 -45289 2 -44911
rect 218 -45022 265 -40668
rect 329 -45022 345 -40668
rect 218 -45038 345 -45022
rect 218 -45162 322 -45038
rect 218 -45178 345 -45162
rect -211 -45290 111 -45289
rect -211 -49420 -210 -45290
rect 110 -49420 111 -45290
rect -211 -49421 111 -49420
rect -102 -49799 2 -49421
rect 218 -49532 265 -45178
rect 329 -49532 345 -45178
rect 218 -49548 345 -49532
rect 218 -49672 322 -49548
rect 218 -49688 345 -49672
rect -211 -49800 111 -49799
rect -211 -53930 -210 -49800
rect 110 -53930 111 -49800
rect -211 -53931 111 -53930
rect -102 -54309 2 -53931
rect 218 -54042 265 -49688
rect 329 -54042 345 -49688
rect 218 -54058 345 -54042
rect 218 -54182 322 -54058
rect 218 -54198 345 -54182
rect -211 -54310 111 -54309
rect -211 -58440 -210 -54310
rect 110 -58440 111 -54310
rect -211 -58441 111 -58440
rect -102 -58819 2 -58441
rect 218 -58552 265 -54198
rect 329 -58552 345 -54198
rect 218 -58568 345 -58552
rect 218 -58692 322 -58568
rect 218 -58708 345 -58692
rect -211 -58820 111 -58819
rect -211 -62950 -210 -58820
rect 110 -62950 111 -58820
rect -211 -62951 111 -62950
rect -102 -63329 2 -62951
rect 218 -63062 265 -58708
rect 329 -63062 345 -58708
rect 218 -63078 345 -63062
rect 218 -63202 322 -63078
rect 218 -63218 345 -63202
rect -211 -63330 111 -63329
rect -211 -67460 -210 -63330
rect 110 -67460 111 -63330
rect -211 -67461 111 -67460
rect -102 -67839 2 -67461
rect 218 -67572 265 -63218
rect 329 -67572 345 -63218
rect 218 -67588 345 -67572
rect 218 -67712 322 -67588
rect 218 -67728 345 -67712
rect -211 -67840 111 -67839
rect -211 -71970 -210 -67840
rect 110 -71970 111 -67840
rect -211 -71971 111 -71970
rect -102 -72349 2 -71971
rect 218 -72082 265 -67728
rect 329 -72082 345 -67728
rect 218 -72098 345 -72082
rect 218 -72222 322 -72098
rect 218 -72238 345 -72222
rect -211 -72350 111 -72349
rect -211 -76480 -210 -72350
rect 110 -76480 111 -72350
rect -211 -76481 111 -76480
rect -102 -76859 2 -76481
rect 218 -76592 265 -72238
rect 329 -76592 345 -72238
rect 218 -76608 345 -76592
rect 218 -76732 322 -76608
rect 218 -76748 345 -76732
rect -211 -76860 111 -76859
rect -211 -80990 -210 -76860
rect 110 -80990 111 -76860
rect -211 -80991 111 -80990
rect -102 -81369 2 -80991
rect 218 -81102 265 -76748
rect 329 -81102 345 -76748
rect 218 -81118 345 -81102
rect 218 -81242 322 -81118
rect 218 -81258 345 -81242
rect -211 -81370 111 -81369
rect -211 -85500 -210 -81370
rect 110 -85500 111 -81370
rect -211 -85501 111 -85500
rect -102 -85879 2 -85501
rect 218 -85612 265 -81258
rect 329 -85612 345 -81258
rect 218 -85628 345 -85612
rect 218 -85752 322 -85628
rect 218 -85768 345 -85752
rect -211 -85880 111 -85879
rect -211 -90010 -210 -85880
rect 110 -90010 111 -85880
rect -211 -90011 111 -90010
rect -102 -90389 2 -90011
rect 218 -90122 265 -85768
rect 329 -90122 345 -85768
rect 218 -90138 345 -90122
rect 218 -90262 322 -90138
rect 218 -90278 345 -90262
rect -211 -90390 111 -90389
rect -211 -94520 -210 -90390
rect 110 -94520 111 -90390
rect -211 -94521 111 -94520
rect -102 -94899 2 -94521
rect 218 -94632 265 -90278
rect 329 -94632 345 -90278
rect 218 -94648 345 -94632
rect 218 -94772 322 -94648
rect 218 -94788 345 -94772
rect -211 -94900 111 -94899
rect -211 -99030 -210 -94900
rect 110 -99030 111 -94900
rect -211 -99031 111 -99030
rect -102 -99409 2 -99031
rect 218 -99142 265 -94788
rect 329 -99142 345 -94788
rect 218 -99158 345 -99142
rect 218 -99282 322 -99158
rect 218 -99298 345 -99282
rect -211 -99410 111 -99409
rect -211 -103540 -210 -99410
rect 110 -103540 111 -99410
rect -211 -103541 111 -103540
rect -102 -103919 2 -103541
rect 218 -103652 265 -99298
rect 329 -103652 345 -99298
rect 218 -103668 345 -103652
rect 218 -103792 322 -103668
rect 218 -103808 345 -103792
rect -211 -103920 111 -103919
rect -211 -108050 -210 -103920
rect 110 -108050 111 -103920
rect -211 -108051 111 -108050
rect -102 -108429 2 -108051
rect 218 -108162 265 -103808
rect 329 -108162 345 -103808
rect 218 -108178 345 -108162
rect 218 -108302 322 -108178
rect 218 -108318 345 -108302
rect -211 -108430 111 -108429
rect -211 -112560 -210 -108430
rect 110 -112560 111 -108430
rect -211 -112561 111 -112560
rect -102 -112939 2 -112561
rect 218 -112672 265 -108318
rect 329 -112672 345 -108318
rect 218 -112688 345 -112672
rect 218 -112812 322 -112688
rect 218 -112828 345 -112812
rect -211 -112940 111 -112939
rect -211 -117070 -210 -112940
rect 110 -117070 111 -112940
rect -211 -117071 111 -117070
rect -102 -117449 2 -117071
rect 218 -117182 265 -112828
rect 329 -117182 345 -112828
rect 218 -117198 345 -117182
rect 218 -117322 322 -117198
rect 218 -117338 345 -117322
rect -211 -117450 111 -117449
rect -211 -121580 -210 -117450
rect 110 -121580 111 -117450
rect -211 -121581 111 -121580
rect -102 -121959 2 -121581
rect 218 -121692 265 -117338
rect 329 -121692 345 -117338
rect 218 -121708 345 -121692
rect 218 -121832 322 -121708
rect 218 -121848 345 -121832
rect -211 -121960 111 -121959
rect -211 -126090 -210 -121960
rect 110 -126090 111 -121960
rect -211 -126091 111 -126090
rect -102 -126469 2 -126091
rect 218 -126202 265 -121848
rect 329 -126202 345 -121848
rect 218 -126218 345 -126202
rect 218 -126342 322 -126218
rect 218 -126358 345 -126342
rect -211 -126470 111 -126469
rect -211 -130600 -210 -126470
rect 110 -130600 111 -126470
rect -211 -130601 111 -130600
rect -102 -130979 2 -130601
rect 218 -130712 265 -126358
rect 329 -130712 345 -126358
rect 218 -130728 345 -130712
rect 218 -130852 322 -130728
rect 218 -130868 345 -130852
rect -211 -130980 111 -130979
rect -211 -135110 -210 -130980
rect 110 -135110 111 -130980
rect -211 -135111 111 -135110
rect -102 -135489 2 -135111
rect 218 -135222 265 -130868
rect 329 -135222 345 -130868
rect 218 -135238 345 -135222
rect 218 -135362 322 -135238
rect 218 -135378 345 -135362
rect -211 -135490 111 -135489
rect -211 -139620 -210 -135490
rect 110 -139620 111 -135490
rect -211 -139621 111 -139620
rect -102 -139999 2 -139621
rect 218 -139732 265 -135378
rect 329 -139732 345 -135378
rect 218 -139748 345 -139732
rect 218 -139872 322 -139748
rect 218 -139888 345 -139872
rect -211 -140000 111 -139999
rect -211 -144130 -210 -140000
rect 110 -144130 111 -140000
rect -211 -144131 111 -144130
rect -102 -144509 2 -144131
rect 218 -144242 265 -139888
rect 329 -144242 345 -139888
rect 218 -144258 345 -144242
rect 218 -144382 322 -144258
rect 218 -144398 345 -144382
rect -211 -144510 111 -144509
rect -211 -148640 -210 -144510
rect 110 -148640 111 -144510
rect -211 -148641 111 -148640
rect -102 -149019 2 -148641
rect 218 -148752 265 -144398
rect 329 -148752 345 -144398
rect 218 -148768 345 -148752
rect 218 -148892 322 -148768
rect 218 -148908 345 -148892
rect -211 -149020 111 -149019
rect -211 -153150 -210 -149020
rect 110 -153150 111 -149020
rect -211 -153151 111 -153150
rect -102 -153529 2 -153151
rect 218 -153262 265 -148908
rect 329 -153262 345 -148908
rect 218 -153278 345 -153262
rect 218 -153402 322 -153278
rect 218 -153418 345 -153402
rect -211 -153530 111 -153529
rect -211 -157660 -210 -153530
rect 110 -157660 111 -153530
rect -211 -157661 111 -157660
rect -102 -158039 2 -157661
rect 218 -157772 265 -153418
rect 329 -157772 345 -153418
rect 218 -157788 345 -157772
rect 218 -157912 322 -157788
rect 218 -157928 345 -157912
rect -211 -158040 111 -158039
rect -211 -162170 -210 -158040
rect 110 -162170 111 -158040
rect -211 -162171 111 -162170
rect -102 -162549 2 -162171
rect 218 -162282 265 -157928
rect 329 -162282 345 -157928
rect 218 -162298 345 -162282
rect 218 -162422 322 -162298
rect 218 -162438 345 -162422
rect -211 -162550 111 -162549
rect -211 -166680 -210 -162550
rect 110 -166680 111 -162550
rect -211 -166681 111 -166680
rect -102 -167059 2 -166681
rect 218 -166792 265 -162438
rect 329 -166792 345 -162438
rect 218 -166808 345 -166792
rect 218 -166932 322 -166808
rect 218 -166948 345 -166932
rect -211 -167060 111 -167059
rect -211 -171190 -210 -167060
rect 110 -171190 111 -167060
rect -211 -171191 111 -171190
rect -102 -171569 2 -171191
rect 218 -171302 265 -166948
rect 329 -171302 345 -166948
rect 218 -171318 345 -171302
rect 218 -171442 322 -171318
rect 218 -171458 345 -171442
rect -211 -171570 111 -171569
rect -211 -175700 -210 -171570
rect 110 -175700 111 -171570
rect -211 -175701 111 -175700
rect -102 -176079 2 -175701
rect 218 -175812 265 -171458
rect 329 -175812 345 -171458
rect 218 -175828 345 -175812
rect 218 -175952 322 -175828
rect 218 -175968 345 -175952
rect -211 -176080 111 -176079
rect -211 -180210 -210 -176080
rect 110 -180210 111 -176080
rect -211 -180211 111 -180210
rect -102 -180589 2 -180211
rect 218 -180322 265 -175968
rect 329 -180322 345 -175968
rect 218 -180338 345 -180322
rect 218 -180462 322 -180338
rect 218 -180478 345 -180462
rect -211 -180590 111 -180589
rect -211 -184720 -210 -180590
rect 110 -184720 111 -180590
rect -211 -184721 111 -184720
rect -102 -185099 2 -184721
rect 218 -184832 265 -180478
rect 329 -184832 345 -180478
rect 218 -184848 345 -184832
rect 218 -184972 322 -184848
rect 218 -184988 345 -184972
rect -211 -185100 111 -185099
rect -211 -189230 -210 -185100
rect 110 -189230 111 -185100
rect -211 -189231 111 -189230
rect -102 -189609 2 -189231
rect 218 -189342 265 -184988
rect 329 -189342 345 -184988
rect 218 -189358 345 -189342
rect 218 -189482 322 -189358
rect 218 -189498 345 -189482
rect -211 -189610 111 -189609
rect -211 -193740 -210 -189610
rect 110 -193740 111 -189610
rect -211 -193741 111 -193740
rect -102 -194119 2 -193741
rect 218 -193852 265 -189498
rect 329 -193852 345 -189498
rect 218 -193868 345 -193852
rect 218 -193992 322 -193868
rect 218 -194008 345 -193992
rect -211 -194120 111 -194119
rect -211 -198250 -210 -194120
rect 110 -198250 111 -194120
rect -211 -198251 111 -198250
rect -102 -198629 2 -198251
rect 218 -198362 265 -194008
rect 329 -198362 345 -194008
rect 218 -198378 345 -198362
rect 218 -198502 322 -198378
rect 218 -198518 345 -198502
rect -211 -198630 111 -198629
rect -211 -202760 -210 -198630
rect 110 -202760 111 -198630
rect -211 -202761 111 -202760
rect -102 -203139 2 -202761
rect 218 -202872 265 -198518
rect 329 -202872 345 -198518
rect 218 -202888 345 -202872
rect 218 -203012 322 -202888
rect 218 -203028 345 -203012
rect -211 -203140 111 -203139
rect -211 -207270 -210 -203140
rect 110 -207270 111 -203140
rect -211 -207271 111 -207270
rect -102 -207649 2 -207271
rect 218 -207382 265 -203028
rect 329 -207382 345 -203028
rect 218 -207398 345 -207382
rect 218 -207522 322 -207398
rect 218 -207538 345 -207522
rect -211 -207650 111 -207649
rect -211 -211780 -210 -207650
rect 110 -211780 111 -207650
rect -211 -211781 111 -211780
rect -102 -212159 2 -211781
rect 218 -211892 265 -207538
rect 329 -211892 345 -207538
rect 218 -211908 345 -211892
rect 218 -212032 322 -211908
rect 218 -212048 345 -212032
rect -211 -212160 111 -212159
rect -211 -216290 -210 -212160
rect 110 -216290 111 -212160
rect -211 -216291 111 -216290
rect -102 -216669 2 -216291
rect 218 -216402 265 -212048
rect 329 -216402 345 -212048
rect 218 -216418 345 -216402
rect 218 -216542 322 -216418
rect 218 -216558 345 -216542
rect -211 -216670 111 -216669
rect -211 -220800 -210 -216670
rect 110 -220800 111 -216670
rect -211 -220801 111 -220800
rect -102 -221179 2 -220801
rect 218 -220912 265 -216558
rect 329 -220912 345 -216558
rect 218 -220928 345 -220912
rect 218 -221052 322 -220928
rect 218 -221068 345 -221052
rect -211 -221180 111 -221179
rect -211 -225310 -210 -221180
rect 110 -225310 111 -221180
rect -211 -225311 111 -225310
rect -102 -225689 2 -225311
rect 218 -225422 265 -221068
rect 329 -225422 345 -221068
rect 218 -225438 345 -225422
rect 218 -225562 322 -225438
rect 218 -225578 345 -225562
rect -211 -225690 111 -225689
rect -211 -229820 -210 -225690
rect 110 -229820 111 -225690
rect -211 -229821 111 -229820
rect -102 -230199 2 -229821
rect 218 -229932 265 -225578
rect 329 -229932 345 -225578
rect 218 -229948 345 -229932
rect 218 -230072 322 -229948
rect 218 -230088 345 -230072
rect -211 -230200 111 -230199
rect -211 -234330 -210 -230200
rect 110 -234330 111 -230200
rect -211 -234331 111 -234330
rect -102 -234709 2 -234331
rect 218 -234442 265 -230088
rect 329 -234442 345 -230088
rect 218 -234458 345 -234442
rect 218 -234582 322 -234458
rect 218 -234598 345 -234582
rect -211 -234710 111 -234709
rect -211 -238840 -210 -234710
rect 110 -238840 111 -234710
rect -211 -238841 111 -238840
rect -102 -239219 2 -238841
rect 218 -238952 265 -234598
rect 329 -238952 345 -234598
rect 218 -238968 345 -238952
rect 218 -239092 322 -238968
rect 218 -239108 345 -239092
rect -211 -239220 111 -239219
rect -211 -243350 -210 -239220
rect 110 -243350 111 -239220
rect -211 -243351 111 -243350
rect -102 -243729 2 -243351
rect 218 -243462 265 -239108
rect 329 -243462 345 -239108
rect 218 -243478 345 -243462
rect 218 -243602 322 -243478
rect 218 -243618 345 -243602
rect -211 -243730 111 -243729
rect -211 -247860 -210 -243730
rect 110 -247860 111 -243730
rect -211 -247861 111 -247860
rect -102 -248239 2 -247861
rect 218 -247972 265 -243618
rect 329 -247972 345 -243618
rect 218 -247988 345 -247972
rect 218 -248112 322 -247988
rect 218 -248128 345 -248112
rect -211 -248240 111 -248239
rect -211 -252370 -210 -248240
rect 110 -252370 111 -248240
rect -211 -252371 111 -252370
rect -102 -252749 2 -252371
rect 218 -252482 265 -248128
rect 329 -252482 345 -248128
rect 218 -252498 345 -252482
rect 218 -252622 322 -252498
rect 218 -252638 345 -252622
rect -211 -252750 111 -252749
rect -211 -256880 -210 -252750
rect 110 -256880 111 -252750
rect -211 -256881 111 -256880
rect -102 -257259 2 -256881
rect 218 -256992 265 -252638
rect 329 -256992 345 -252638
rect 218 -257008 345 -256992
rect 218 -257132 322 -257008
rect 218 -257148 345 -257132
rect -211 -257260 111 -257259
rect -211 -261390 -210 -257260
rect 110 -261390 111 -257260
rect -211 -261391 111 -261390
rect -102 -261769 2 -261391
rect 218 -261502 265 -257148
rect 329 -261502 345 -257148
rect 218 -261518 345 -261502
rect 218 -261642 322 -261518
rect 218 -261658 345 -261642
rect -211 -261770 111 -261769
rect -211 -265900 -210 -261770
rect 110 -265900 111 -261770
rect -211 -265901 111 -265900
rect -102 -266279 2 -265901
rect 218 -266012 265 -261658
rect 329 -266012 345 -261658
rect 218 -266028 345 -266012
rect 218 -266152 322 -266028
rect 218 -266168 345 -266152
rect -211 -266280 111 -266279
rect -211 -270410 -210 -266280
rect 110 -270410 111 -266280
rect -211 -270411 111 -270410
rect -102 -270789 2 -270411
rect 218 -270522 265 -266168
rect 329 -270522 345 -266168
rect 218 -270538 345 -270522
rect 218 -270662 322 -270538
rect 218 -270678 345 -270662
rect -211 -270790 111 -270789
rect -211 -274920 -210 -270790
rect 110 -274920 111 -270790
rect -211 -274921 111 -274920
rect -102 -275299 2 -274921
rect 218 -275032 265 -270678
rect 329 -275032 345 -270678
rect 218 -275048 345 -275032
rect 218 -275172 322 -275048
rect 218 -275188 345 -275172
rect -211 -275300 111 -275299
rect -211 -279430 -210 -275300
rect 110 -279430 111 -275300
rect -211 -279431 111 -279430
rect -102 -279809 2 -279431
rect 218 -279542 265 -275188
rect 329 -279542 345 -275188
rect 218 -279558 345 -279542
rect 218 -279682 322 -279558
rect 218 -279698 345 -279682
rect -211 -279810 111 -279809
rect -211 -283940 -210 -279810
rect 110 -283940 111 -279810
rect -211 -283941 111 -283940
rect -102 -284319 2 -283941
rect 218 -284052 265 -279698
rect 329 -284052 345 -279698
rect 218 -284068 345 -284052
rect 218 -284192 322 -284068
rect 218 -284208 345 -284192
rect -211 -284320 111 -284319
rect -211 -288450 -210 -284320
rect 110 -288450 111 -284320
rect -211 -288451 111 -288450
rect -102 -288640 2 -288451
rect 218 -288562 265 -284208
rect 329 -288562 345 -284208
rect 218 -288578 345 -288562
rect 218 -288640 322 -288578
<< properties >>
string FIXED_BBOX -350 284180 250 288590
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 128 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
