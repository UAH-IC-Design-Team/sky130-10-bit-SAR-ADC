magic
tech sky130A
magscale 1 2
timestamp 1668208340
<< nwell >>
rect 4690 -3340 5180 -2700
rect 8370 -3340 8860 -2700
rect 5020 -4620 5550 -3640
rect 8000 -4620 8530 -3640
<< psubdiff >>
rect 4410 -2630 4510 -2606
rect 4410 -2894 4510 -2870
rect 9040 -2610 9140 -2586
rect 9040 -2874 9140 -2850
rect 4410 -4680 4510 -4656
rect 4410 -4944 4510 -4920
rect 9040 -4690 9140 -4666
rect 9040 -4954 9140 -4930
<< nsubdiff >>
rect 4820 -3070 4850 -2970
rect 4980 -3070 5010 -2970
rect 8540 -3070 8570 -2970
rect 8700 -3070 8730 -2970
rect 5080 -4380 5110 -4300
rect 5320 -4380 5350 -4300
rect 8200 -4380 8230 -4300
rect 8440 -4380 8470 -4300
<< psubdiffcont >>
rect 4410 -2870 4510 -2630
rect 9040 -2850 9140 -2610
rect 4410 -4920 4510 -4680
rect 9040 -4930 9140 -4690
<< nsubdiffcont >>
rect 4850 -3070 4980 -2970
rect 8570 -3070 8700 -2970
rect 5110 -4380 5320 -4300
rect 8230 -4380 8440 -4300
<< locali >>
rect 9040 -2610 9140 -2594
rect 4410 -2630 4510 -2614
rect 9040 -2866 9140 -2850
rect 4410 -2886 4510 -2870
rect 4830 -3070 4850 -2970
rect 4980 -3070 5000 -2970
rect 8550 -3070 8570 -2970
rect 8700 -3070 8720 -2970
rect 5090 -4380 5110 -4300
rect 5320 -4380 5340 -4300
rect 8210 -4380 8230 -4300
rect 8440 -4380 8460 -4300
rect 4410 -4680 4510 -4664
rect 4410 -4936 4510 -4920
rect 9040 -4690 9140 -4674
rect 9040 -4946 9140 -4930
<< viali >>
rect 4420 -2870 4500 -2630
rect 9050 -2850 9130 -2610
rect 4850 -3070 4980 -2970
rect 8570 -3070 8700 -2970
rect 5130 -4370 5300 -4310
rect 8250 -4370 8420 -4310
rect 4420 -4920 4500 -4680
rect 9050 -4930 9130 -4690
<< metal1 >>
rect 4670 -2320 4850 -2310
rect 4670 -2390 4680 -2320
rect 4750 -2390 4770 -2320
rect 4840 -2390 4850 -2320
rect 4670 -2400 4850 -2390
rect 8700 -2320 8880 -2310
rect 8700 -2390 8710 -2320
rect 8780 -2390 8800 -2320
rect 8870 -2390 8880 -2320
rect 8700 -2400 8880 -2390
rect 4360 -2450 4510 -2440
rect 4420 -2550 4450 -2450
rect 4360 -2630 4510 -2550
rect 4360 -2870 4420 -2630
rect 4500 -2870 4510 -2630
rect 4360 -4680 4510 -2870
rect 4560 -2650 4640 -2640
rect 4612 -2710 4640 -2650
rect 4560 -2730 4640 -2710
rect 4612 -2790 4640 -2730
rect 4560 -3630 4640 -2790
rect 4680 -3530 4750 -2400
rect 5650 -2450 5820 -2440
rect 4780 -2470 4960 -2460
rect 4780 -2530 4790 -2470
rect 4950 -2530 4960 -2470
rect 4780 -2540 4960 -2530
rect 5650 -2530 5670 -2450
rect 5730 -2530 5750 -2450
rect 5810 -2530 5820 -2450
rect 5650 -2560 5820 -2530
rect 4800 -2650 4940 -2580
rect 4930 -2660 4940 -2650
rect 4930 -2710 5690 -2660
rect 4800 -2790 4940 -2710
rect 4820 -2960 5030 -2830
rect 5150 -2960 5470 -2910
rect 5620 -2950 5690 -2710
rect 4820 -2970 5230 -2960
rect 4820 -3080 4830 -2970
rect 5010 -3080 5040 -2970
rect 5220 -3080 5230 -2970
rect 5740 -2980 5820 -2560
rect 5360 -3050 5630 -2990
rect 5360 -3070 5420 -3050
rect 5680 -3070 5820 -2980
rect 7720 -2450 7900 -2440
rect 7720 -2530 7730 -2450
rect 7800 -2530 7820 -2450
rect 7890 -2530 7900 -2450
rect 7720 -2560 7900 -2530
rect 8590 -2470 8770 -2460
rect 8590 -2530 8600 -2470
rect 8760 -2530 8770 -2470
rect 8590 -2540 8770 -2530
rect 7720 -2980 7810 -2560
rect 8610 -2650 8750 -2580
rect 8610 -2660 8620 -2650
rect 7860 -2710 8620 -2660
rect 7860 -2950 7930 -2710
rect 8610 -2790 8750 -2710
rect 8080 -2960 8400 -2910
rect 8520 -2960 8730 -2830
rect 8320 -2970 8730 -2960
rect 7720 -3060 7870 -2980
rect 7920 -3050 8190 -2990
rect 8130 -3070 8190 -3050
rect 4820 -3100 5230 -3080
rect 4820 -3210 5030 -3100
rect 4790 -3350 4960 -3260
rect 4790 -3420 5080 -3350
rect 4790 -3480 4960 -3420
rect 4560 -3710 4720 -3630
rect 4360 -4920 4420 -4680
rect 4500 -4920 4510 -4680
rect 4650 -4910 4720 -3710
rect 4860 -3810 4960 -3520
rect 4820 -3820 4960 -3810
rect 4820 -3890 4830 -3820
rect 4940 -3890 4960 -3820
rect 4820 -3930 4960 -3890
rect 4820 -4000 4830 -3930
rect 4940 -4000 4960 -3930
rect 4820 -4010 4960 -4000
rect 4360 -4960 4510 -4920
rect 4750 -4960 4820 -4210
rect 4360 -5070 4820 -4960
rect 4860 -4960 4960 -4010
rect 5010 -4470 5080 -3420
rect 5150 -3660 5230 -3100
rect 8320 -3080 8330 -2970
rect 8510 -3080 8540 -2970
rect 8720 -3080 8730 -2970
rect 8320 -3100 8730 -3080
rect 5270 -3180 5520 -3110
rect 5450 -3240 5520 -3180
rect 8030 -3180 8280 -3110
rect 8030 -3240 8100 -3180
rect 5450 -3310 5650 -3240
rect 5120 -3730 5230 -3660
rect 5580 -3730 5650 -3310
rect 5120 -4120 5190 -3730
rect 5360 -3780 5650 -3730
rect 5242 -4210 5320 -3790
rect 5220 -4230 5320 -4210
rect 5110 -4240 5320 -4230
rect 5110 -4310 5120 -4240
rect 5310 -4310 5320 -4240
rect 5110 -4350 5130 -4310
rect 5300 -4350 5320 -4310
rect 5110 -4420 5120 -4350
rect 5310 -4420 5320 -4350
rect 5110 -4430 5320 -4420
rect 5010 -4560 5130 -4470
rect 5050 -4750 5130 -4560
rect 5180 -4580 5320 -4430
rect 5360 -4000 5420 -3780
rect 5580 -4000 5650 -3780
rect 5360 -4050 5650 -4000
rect 5360 -4170 5420 -4050
rect 5580 -4170 5650 -4050
rect 5360 -4220 5650 -4170
rect 5360 -4440 5420 -4220
rect 5580 -4440 5650 -4220
rect 5360 -4490 5650 -4440
rect 5580 -4650 5650 -4490
rect 5270 -4710 5650 -4650
rect 5050 -4840 5280 -4750
rect 5330 -4960 5480 -4740
rect 5690 -4750 6060 -3240
rect 5520 -4890 6060 -4750
rect 6180 -4890 6570 -3240
rect 6980 -4890 7370 -3240
rect 7490 -4750 7860 -3240
rect 7900 -3310 8100 -3240
rect 7900 -3730 7970 -3310
rect 8320 -3660 8400 -3100
rect 8520 -3210 8730 -3100
rect 8590 -3350 8760 -3260
rect 8470 -3420 8760 -3350
rect 8320 -3730 8430 -3660
rect 7900 -3780 8190 -3730
rect 7900 -4000 7970 -3780
rect 8130 -4000 8190 -3780
rect 7900 -4050 8190 -4000
rect 7900 -4170 7970 -4050
rect 8130 -4170 8190 -4050
rect 7900 -4220 8190 -4170
rect 7900 -4440 7970 -4220
rect 8130 -4440 8190 -4220
rect 7900 -4490 8190 -4440
rect 8230 -4210 8308 -3790
rect 8360 -4120 8430 -3730
rect 8230 -4230 8330 -4210
rect 8230 -4240 8440 -4230
rect 8230 -4310 8240 -4240
rect 8430 -4310 8440 -4240
rect 8230 -4350 8250 -4310
rect 8420 -4350 8440 -4310
rect 8230 -4420 8240 -4350
rect 8430 -4420 8440 -4350
rect 8230 -4430 8440 -4420
rect 7900 -4650 7970 -4490
rect 8230 -4580 8370 -4430
rect 8470 -4470 8540 -3420
rect 8590 -3480 8760 -3420
rect 8420 -4560 8540 -4470
rect 8590 -3810 8690 -3520
rect 8800 -3530 8870 -2400
rect 9040 -2450 9190 -2440
rect 9100 -2550 9130 -2450
rect 9040 -2610 9190 -2550
rect 8910 -2650 8990 -2640
rect 8910 -2710 8938 -2650
rect 8910 -2730 8990 -2710
rect 8910 -2790 8938 -2730
rect 8910 -3630 8990 -2790
rect 8830 -3710 8990 -3630
rect 9040 -2850 9050 -2610
rect 9130 -2850 9190 -2610
rect 8590 -3820 8730 -3810
rect 8590 -3890 8600 -3820
rect 8720 -3890 8730 -3820
rect 8590 -3930 8730 -3890
rect 8590 -4000 8600 -3930
rect 8720 -4000 8730 -3930
rect 8590 -4010 8730 -4000
rect 7900 -4710 8280 -4650
rect 7490 -4890 8030 -4750
rect 4860 -5070 5480 -4960
rect 8070 -4960 8220 -4740
rect 8420 -4750 8500 -4560
rect 8270 -4840 8500 -4750
rect 8590 -4960 8690 -4010
rect 8070 -5070 8690 -4960
rect 8730 -4960 8800 -4210
rect 8830 -4910 8900 -3710
rect 9040 -4690 9190 -2850
rect 9040 -4930 9050 -4690
rect 9130 -4930 9190 -4690
rect 9040 -4960 9190 -4930
rect 8730 -5070 9190 -4960
<< via1 >>
rect 4680 -2390 4750 -2320
rect 4770 -2390 4840 -2320
rect 8710 -2390 8780 -2320
rect 8800 -2390 8870 -2320
rect 4360 -2550 4420 -2450
rect 4450 -2550 4510 -2450
rect 4560 -2710 4612 -2650
rect 4560 -2790 4612 -2730
rect 4790 -2530 4950 -2470
rect 5670 -2530 5730 -2450
rect 5750 -2530 5810 -2450
rect 4800 -2710 4930 -2650
rect 4830 -3070 4850 -2970
rect 4850 -3070 4980 -2970
rect 4980 -3070 5010 -2970
rect 4830 -3080 5010 -3070
rect 5040 -3080 5220 -2970
rect 7730 -2530 7800 -2450
rect 7820 -2530 7890 -2450
rect 8600 -2530 8760 -2470
rect 8620 -2710 8750 -2650
rect 4830 -3890 4940 -3820
rect 4830 -4000 4940 -3930
rect 8330 -3080 8510 -2970
rect 8540 -3070 8570 -2970
rect 8570 -3070 8700 -2970
rect 8700 -3070 8720 -2970
rect 8540 -3080 8720 -3070
rect 5120 -4310 5310 -4240
rect 5120 -4370 5130 -4350
rect 5130 -4370 5300 -4350
rect 5300 -4370 5310 -4350
rect 5120 -4420 5310 -4370
rect 8240 -4310 8430 -4240
rect 8240 -4370 8250 -4350
rect 8250 -4370 8420 -4350
rect 8420 -4370 8430 -4350
rect 8240 -4420 8430 -4370
rect 9040 -2550 9100 -2450
rect 9130 -2550 9190 -2450
rect 8938 -2710 8990 -2650
rect 8938 -2790 8990 -2730
rect 8600 -3890 8720 -3820
rect 8600 -4000 8720 -3930
<< metal2 >>
rect 4670 -2320 8880 -2310
rect 4670 -2390 4680 -2320
rect 4750 -2390 4770 -2320
rect 4840 -2390 8710 -2320
rect 8780 -2390 8800 -2320
rect 8870 -2390 8880 -2320
rect 4670 -2400 8880 -2390
rect 4360 -2450 9190 -2440
rect 4420 -2550 4450 -2450
rect 4510 -2470 5670 -2450
rect 4510 -2530 4790 -2470
rect 4950 -2530 5670 -2470
rect 5730 -2530 5750 -2450
rect 5810 -2530 7730 -2450
rect 7800 -2530 7820 -2450
rect 7890 -2470 9040 -2450
rect 7890 -2530 8600 -2470
rect 8760 -2530 9040 -2470
rect 4510 -2550 9040 -2530
rect 9100 -2550 9130 -2450
rect 4360 -2560 9190 -2550
rect 4550 -2650 4940 -2640
rect 4550 -2710 4560 -2650
rect 4612 -2710 4800 -2650
rect 4930 -2710 4940 -2650
rect 4550 -2720 4940 -2710
rect 8610 -2650 9000 -2640
rect 8610 -2710 8620 -2650
rect 8750 -2710 8938 -2650
rect 8990 -2710 9000 -2650
rect 8610 -2720 9000 -2710
rect 4550 -2730 4620 -2720
rect 4550 -2790 4560 -2730
rect 4612 -2790 4620 -2730
rect 4550 -2800 4620 -2790
rect 8930 -2730 9000 -2720
rect 8930 -2790 8938 -2730
rect 8990 -2790 9000 -2730
rect 8930 -2800 9000 -2790
rect 4820 -2970 8730 -2960
rect 4820 -3080 4830 -2970
rect 5010 -3080 5040 -2970
rect 5220 -3080 8330 -2970
rect 8510 -3080 8540 -2970
rect 8720 -3080 8730 -2970
rect 4820 -3100 8730 -3080
rect 4330 -3820 4960 -3810
rect 4330 -3890 4340 -3820
rect 4480 -3890 4830 -3820
rect 4940 -3890 4960 -3820
rect 4330 -3930 4960 -3890
rect 4330 -4000 4340 -3930
rect 4480 -4000 4830 -3930
rect 4940 -4000 4960 -3930
rect 4330 -4010 4960 -4000
rect 8590 -3820 9220 -3810
rect 8590 -3890 8600 -3820
rect 8720 -3890 9070 -3820
rect 9210 -3890 9220 -3820
rect 8590 -3930 9220 -3890
rect 8590 -4000 8600 -3930
rect 8720 -4000 9070 -3930
rect 9210 -4000 9220 -3930
rect 8590 -4010 9220 -4000
rect 3990 -4240 5320 -4230
rect 3990 -4310 4010 -4240
rect 4190 -4310 5120 -4240
rect 5310 -4310 5320 -4240
rect 3990 -4340 5320 -4310
rect 3990 -4420 4010 -4340
rect 4190 -4350 5320 -4340
rect 4190 -4420 5120 -4350
rect 5310 -4420 5320 -4350
rect 3990 -4430 5320 -4420
rect 8230 -4240 9560 -4230
rect 8230 -4310 8240 -4240
rect 8430 -4310 9360 -4240
rect 9550 -4310 9560 -4240
rect 8230 -4350 9560 -4310
rect 8230 -4420 8240 -4350
rect 8430 -4420 9360 -4350
rect 9550 -4420 9560 -4350
rect 8230 -4430 9560 -4420
<< via2 >>
rect 4340 -3890 4480 -3820
rect 4340 -4000 4480 -3930
rect 9070 -3890 9210 -3820
rect 9070 -4000 9210 -3930
rect 4010 -4310 4190 -4240
rect 4010 -4420 4190 -4340
rect 9360 -4310 9550 -4240
rect 9360 -4420 9550 -4350
<< metal3 >>
rect -3600 500 4200 900
rect -3600 -1900 -3400 500
rect 4000 -1900 4200 500
rect -3600 -2300 4200 -1900
rect -3600 -4700 -3400 -2300
rect 4000 -4240 4200 -2300
rect 9350 500 17150 900
rect 9350 -1900 9550 500
rect 16950 -1900 17150 500
rect 9350 -2300 17150 -1900
rect 4330 -3820 4490 -3810
rect 4330 -3890 4340 -3820
rect 4480 -3890 4490 -3820
rect 4330 -3930 4490 -3890
rect 4330 -4000 4340 -3930
rect 4480 -4000 4490 -3930
rect 4330 -4010 4490 -4000
rect 9060 -3820 9220 -3810
rect 9060 -3890 9070 -3820
rect 9210 -3890 9220 -3820
rect 9060 -3930 9220 -3890
rect 9060 -4000 9070 -3930
rect 9210 -4000 9220 -3930
rect 9060 -4010 9220 -4000
rect 4000 -4310 4010 -4240
rect 4190 -4310 4200 -4240
rect 4000 -4340 4200 -4310
rect 4000 -4420 4010 -4340
rect 4190 -4420 4200 -4340
rect 4000 -4700 4200 -4420
rect -3600 -5100 4200 -4700
rect 9350 -4240 9550 -2300
rect 9350 -4310 9360 -4240
rect 9350 -4350 9550 -4310
rect 9350 -4420 9360 -4350
rect 9350 -4700 9550 -4420
rect 16950 -4700 17150 -2300
rect 9350 -5100 17150 -4700
<< via3 >>
rect 4340 -3890 4480 -3820
rect 4340 -4000 4480 -3930
rect 9070 -3890 9210 -3820
rect 9070 -4000 9210 -3930
<< metal4 >>
rect -3600 1800 4200 2200
rect -3600 -600 -3400 1800
rect 4000 -600 4200 1800
rect -3600 -1000 4200 -600
rect -3600 -3400 -3400 -1000
rect 4000 -3400 4200 -1000
rect -3600 -3800 4200 -3400
rect 4000 -3810 4200 -3800
rect 9350 1800 17150 2200
rect 9350 -600 9550 1800
rect 16950 -600 17150 1800
rect 9350 -1000 17150 -600
rect 9350 -3400 9550 -1000
rect 16950 -3400 17150 -1000
rect 9350 -3800 17150 -3400
rect 9350 -3810 9550 -3800
rect 4000 -3820 4490 -3810
rect 4000 -3890 4340 -3820
rect 4480 -3890 4490 -3820
rect 4000 -3930 4490 -3890
rect 4000 -4000 4340 -3930
rect 4480 -4000 4490 -3930
rect 4000 -4010 4490 -4000
rect 9060 -3820 9550 -3810
rect 9060 -3890 9070 -3820
rect 9210 -3890 9550 -3820
rect 9060 -3930 9550 -3890
rect 9060 -4000 9070 -3930
rect 9210 -4000 9550 -3930
rect 9060 -4010 9550 -4000
use sky130_fd_pr__nfet_01v8_MRUJZ4  XM1
timestamp 1666807509
transform 0 1 4839 -1 0 -4527
box -413 -179 413 121
use sky130_fd_pr__pfet_01v8_E9NJWS  XM2
timestamp 1666806685
transform 0 1 4915 1 0 -3231
box -109 -225 109 259
use sky130_fd_pr__pfet_01v8_SKSN8V  XM5
timestamp 1666652569
transform 0 -1 5291 -1 0 -4511
box -109 -259 109 225
use sky130_fd_pr__nfet_01v8_P7BBP7  XM8
timestamp 1666651368
transform 0 1 6126 -1 0 -3998
box -749 -543 749 484
use sky130_fd_pr__nfet_01v8_ZWFJZ8  XM9
timestamp 1666724365
transform -1 0 5385 0 -1 -3079
box -125 -179 125 121
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_0
array 0 2 2800 0 2 2600
timestamp 1666650350
transform 0 1 -2300 -1 0 1650
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_1
array 0 2 2800 0 2 2600
timestamp 1666650350
transform 0 -1 15850 -1 0 1650
box -1150 -1100 1149 1100
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_0
timestamp 1666651042
transform -1 0 5503 0 -1 -4802
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_1
timestamp 1666651042
transform 0 1 4838 -1 0 -3497
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_2
timestamp 1666651042
transform 0 1 4838 -1 0 -2557
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_3
timestamp 1666651042
transform 0 -1 8712 -1 0 -2557
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_4
timestamp 1666651042
transform 1 0 8047 0 -1 -4802
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_5
timestamp 1666651042
transform 0 -1 8712 -1 0 -3497
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CME3F  sky130_fd_pr__nfet_01v8_9CME3F_0
timestamp 1666651042
transform 1 0 5303 0 1 -4802
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CME3F  sky130_fd_pr__nfet_01v8_9CME3F_1
timestamp 1666651042
transform 1 0 5653 0 1 -3042
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CME3F  sky130_fd_pr__nfet_01v8_9CME3F_2
timestamp 1666651042
transform -1 0 7897 0 1 -3042
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_9CME3F  sky130_fd_pr__nfet_01v8_9CME3F_3
timestamp 1666651042
transform -1 0 8247 0 1 -4802
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_MRUJZ4  sky130_fd_pr__nfet_01v8_MRUJZ4_0
timestamp 1666807509
transform 0 -1 8711 -1 0 -4527
box -413 -179 413 121
use sky130_fd_pr__nfet_01v8_P7BBP7  sky130_fd_pr__nfet_01v8_P7BBP7_0
timestamp 1666651368
transform 0 -1 7424 -1 0 -3998
box -749 -543 749 484
use sky130_fd_pr__nfet_01v8_ZWFJZ8  sky130_fd_pr__nfet_01v8_ZWFJZ8_0
timestamp 1666724365
transform 1 0 8165 0 -1 -3079
box -125 -179 125 121
use sky130_fd_pr__pfet_01v8_E9NJWS  sky130_fd_pr__pfet_01v8_E9NJWS_0
timestamp 1666806685
transform 0 1 4915 -1 0 -2811
box -109 -225 109 259
use sky130_fd_pr__pfet_01v8_E9NJWS  sky130_fd_pr__pfet_01v8_E9NJWS_1
timestamp 1666806685
transform 0 -1 8635 -1 0 -2811
box -109 -225 109 259
use sky130_fd_pr__pfet_01v8_E9NJWS  sky130_fd_pr__pfet_01v8_E9NJWS_2
timestamp 1666806685
transform 0 -1 8635 1 0 -3231
box -109 -225 109 259
use sky130_fd_pr__pfet_01v8_RQ978N  sky130_fd_pr__pfet_01v8_RQ978N_0
timestamp 1666652569
transform 0 -1 5220 -1 0 -3955
box -305 -200 305 160
use sky130_fd_pr__pfet_01v8_RQ978N  sky130_fd_pr__pfet_01v8_RQ978N_1
timestamp 1666652569
transform 0 1 8330 -1 0 -3955
box -305 -200 305 160
use sky130_fd_pr__pfet_01v8_SKSN8V  sky130_fd_pr__pfet_01v8_SKSN8V_0
timestamp 1666652569
transform 0 1 8259 -1 0 -4511
box -109 -259 109 225
<< labels >>
rlabel metal2 5220 -3100 8330 -2960 1 VDD
port 1 n
rlabel metal1 7490 -4890 7860 -3240 1 Vin_p
port 2 n
rlabel metal1 6980 -4890 7370 -3240 1 Vout_p
port 3 n
rlabel metal2 4950 -2540 8600 -2440 1 VSS
port 4 n
rlabel metal1 6180 -4890 6570 -3240 1 Vout_n
port 5 n
rlabel metal1 5690 -4890 6060 -3240 1 Vin_n
port 6 n
rlabel metal2 4750 -2400 8800 -2310 1 Clk
port 7 n
<< end >>
