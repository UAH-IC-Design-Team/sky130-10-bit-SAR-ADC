magic
tech sky130A
timestamp 1666485801
<< metal4 >>
rect 100 19050 7650 19200
rect 100 19000 150 19050
rect 600 19000 650 19050
rect 1100 19000 1150 19050
rect 1600 19000 1650 19050
rect 2100 19000 2150 19050
rect 2600 19000 2650 19050
rect 3100 19000 3150 19050
rect 3600 19000 3650 19050
rect 4100 19000 4150 19050
rect 4600 19000 4650 19050
rect 5100 19000 5150 19050
rect 5600 19000 5650 19050
rect 6100 19000 6150 19050
rect 6600 19000 6650 19050
rect 7100 19000 7150 19050
rect 7600 19000 7650 19050
rect 8300 19050 11850 19200
rect 8300 19000 8350 19050
rect 8800 19000 8850 19050
rect 9300 19000 9350 19050
rect 9800 19000 9850 19050
rect 10300 19000 10350 19050
rect 10800 19000 10850 19050
rect 11300 19000 11350 19050
rect 11800 19000 11850 19050
rect 12500 19050 20050 19200
rect 12500 19000 12550 19050
rect 13000 19000 13050 19050
rect 13500 19000 13550 19050
rect 14000 19000 14050 19050
rect 14500 19000 14550 19050
rect 15000 19000 15050 19050
rect 15500 19000 15550 19050
rect 16000 19000 16050 19050
rect 16500 19000 16550 19050
rect 17000 19000 17050 19050
rect 17500 19000 17550 19050
rect 18000 19000 18050 19050
rect 18500 19000 18550 19050
rect 19000 19000 19050 19050
rect 19500 19000 19550 19050
rect 20000 19000 20050 19050
rect 20700 19050 24250 19200
rect 20700 19000 20750 19050
rect 21200 19000 21250 19050
rect 21700 19000 21750 19050
rect 22200 19000 22250 19050
rect 22700 19000 22750 19050
rect 23200 19000 23250 19050
rect 23700 19000 23750 19050
rect 24200 19000 24250 19050
rect 24900 19050 26450 19200
rect 24900 19000 24950 19050
rect 25400 19000 25450 19050
rect 25900 19000 25950 19050
rect 26400 19000 26450 19050
rect 27100 19050 27650 19200
rect 27100 19000 27150 19050
rect 27600 19000 27650 19050
rect 28300 19000 28350 19200
rect 29000 19050 30550 19200
rect 29000 19000 29050 19050
rect 29500 19000 29550 19050
rect 30000 19000 30050 19050
rect 30500 19000 30550 19050
rect 31200 19050 31750 19200
rect 31200 19000 31250 19050
rect 31700 19000 31750 19050
rect 32400 19000 32450 19200
rect 33100 2250 34650 2400
rect 35300 2250 35850 2400
rect 36500 2250 36550 2400
rect 37200 2250 38750 2400
rect 39400 2250 39950 2400
rect 40600 2250 40650 2400
rect 41300 2250 41350 2400
rect 300 -50 350 0
rect 800 -50 850 0
rect 1300 -50 1350 0
rect 1800 -50 1850 0
rect 2300 -50 2350 0
rect 2800 -50 2850 0
rect 3300 -50 3350 0
rect 3800 -50 3850 0
rect 4300 -50 4350 0
rect 4800 -50 4850 0
rect 5300 -50 5350 0
rect 5800 -50 5850 0
rect 6300 -50 6350 0
rect 6800 -50 6850 0
rect 7300 -50 7350 0
rect 7800 -50 7850 0
rect 8500 -50 8550 0
rect 9000 -50 9050 0
rect 9500 -50 9550 0
rect 10000 -50 10050 0
rect 10500 -50 10550 0
rect 11000 -50 11050 0
rect 11500 -50 11550 0
rect 12000 -50 12050 0
rect 12700 -50 12750 0
rect 13200 -50 13250 0
rect 13700 -50 13750 0
rect 14200 -50 14250 0
rect 14700 -50 14750 0
rect 15200 -50 15250 0
rect 15700 -50 15750 0
rect 16200 -50 16250 0
rect 16700 -50 16750 0
rect 17200 -50 17250 0
rect 17700 -50 17750 0
rect 18200 -50 18250 0
rect 18700 -50 18750 0
rect 19200 -50 19250 0
rect 19700 -50 19750 0
rect 20200 -50 20250 0
rect 20900 -50 20950 0
rect 21400 -50 21450 0
rect 21900 -50 21950 0
rect 22400 -50 22450 0
rect 22900 -50 22950 0
rect 23400 -50 23450 0
rect 23900 -50 23950 0
rect 24400 -50 24450 0
rect 25100 -50 25150 0
rect 25600 -50 25650 0
rect 26100 -50 26150 0
rect 26600 -50 26650 0
rect 27300 -50 27350 0
rect 27800 -50 27850 0
rect 28500 -50 28550 0
rect 29200 -50 29250 0
rect 29700 -50 29750 0
rect 30200 -50 30250 0
rect 30700 -50 30750 0
rect 31400 -50 31450 0
rect 31900 -50 31950 0
rect 32600 -50 32650 0
rect 33300 -50 33350 0
rect 33800 -50 33850 0
rect 34300 -50 34350 0
rect 34800 -50 34850 0
rect 35500 -50 35550 0
rect 36000 -50 36050 0
rect 36700 -50 36750 0
rect 37400 -50 37450 0
rect 37900 -50 37950 0
rect 38400 -50 38450 0
rect 38900 -50 38950 0
rect 39600 -50 39650 0
rect 40100 -50 40150 0
rect 40800 -50 40850 0
rect 41500 -50 41550 0
rect 300 -200 41550 -50
rect 300 -950 41550 -800
rect 300 -1000 350 -950
rect 800 -1000 850 -950
rect 1300 -1000 1350 -950
rect 1800 -1000 1850 -950
rect 2300 -1000 2350 -950
rect 2800 -1000 2850 -950
rect 3300 -1000 3350 -950
rect 3800 -1000 3850 -950
rect 4300 -1000 4350 -950
rect 4800 -1000 4850 -950
rect 5300 -1000 5350 -950
rect 5800 -1000 5850 -950
rect 6300 -1000 6350 -950
rect 6800 -1000 6850 -950
rect 7300 -1000 7350 -950
rect 7800 -1000 7850 -950
rect 8500 -1000 8550 -950
rect 9000 -1000 9050 -950
rect 9500 -1000 9550 -950
rect 10000 -1000 10050 -950
rect 10500 -1000 10550 -950
rect 11000 -1000 11050 -950
rect 11500 -1000 11550 -950
rect 12000 -1000 12050 -950
rect 12700 -1000 12750 -950
rect 13200 -1000 13250 -950
rect 13700 -1000 13750 -950
rect 14200 -1000 14250 -950
rect 14700 -1000 14750 -950
rect 15200 -1000 15250 -950
rect 15700 -1000 15750 -950
rect 16200 -1000 16250 -950
rect 16700 -1000 16750 -950
rect 17200 -1000 17250 -950
rect 17700 -1000 17750 -950
rect 18200 -1000 18250 -950
rect 18700 -1000 18750 -950
rect 19200 -1000 19250 -950
rect 19700 -1000 19750 -950
rect 20200 -1000 20250 -950
rect 20900 -1000 20950 -950
rect 21400 -1000 21450 -950
rect 21900 -1000 21950 -950
rect 22400 -1000 22450 -950
rect 22900 -1000 22950 -950
rect 23400 -1000 23450 -950
rect 23900 -1000 23950 -950
rect 24400 -1000 24450 -950
rect 25100 -1000 25150 -950
rect 25600 -1000 25650 -950
rect 26100 -1000 26150 -950
rect 26600 -1000 26650 -950
rect 27300 -1000 27350 -950
rect 27800 -1000 27850 -950
rect 28500 -1000 28550 -950
rect 29200 -1000 29250 -950
rect 29700 -1000 29750 -950
rect 30200 -1000 30250 -950
rect 30700 -1000 30750 -950
rect 31400 -1000 31450 -950
rect 31900 -1000 31950 -950
rect 32600 -1000 32650 -950
rect 33300 -1000 33350 -950
rect 33800 -1000 33850 -950
rect 34300 -1000 34350 -950
rect 34800 -1000 34850 -950
rect 35500 -1000 35550 -950
rect 36000 -1000 36050 -950
rect 36700 -1000 36750 -950
rect 37400 -1000 37450 -950
rect 37900 -1000 37950 -950
rect 38400 -1000 38450 -950
rect 38900 -1000 38950 -950
rect 39600 -1000 39650 -950
rect 40100 -1000 40150 -950
rect 40800 -1000 40850 -950
rect 41500 -1000 41550 -950
rect 33100 -3395 34650 -3245
rect 35300 -3395 35850 -3245
rect 36500 -3395 36550 -3245
rect 37200 -3395 38750 -3245
rect 39400 -3395 39950 -3245
rect 40600 -3395 40650 -3245
rect 41300 -3395 41350 -3245
rect 100 -20050 150 -19950
rect 600 -20050 650 -19950
rect 1100 -20050 1150 -19950
rect 1600 -20050 1650 -19950
rect 2100 -20050 2150 -19950
rect 2600 -20050 2650 -19950
rect 3100 -20050 3150 -19950
rect 3600 -20050 3650 -19950
rect 4100 -20050 4150 -19950
rect 4600 -20050 4650 -19950
rect 5100 -20050 5150 -19950
rect 5600 -20050 5650 -19950
rect 6100 -20050 6150 -19950
rect 6600 -20050 6650 -19950
rect 7100 -20050 7150 -19950
rect 7600 -20050 7650 -19950
rect 100 -20200 7650 -20050
rect 8300 -20050 8350 -19950
rect 8800 -20050 8850 -19950
rect 9300 -20050 9350 -19950
rect 9800 -20050 9850 -19950
rect 10300 -20050 10350 -19950
rect 10800 -20050 10850 -19950
rect 11300 -20050 11350 -19950
rect 11800 -20050 11850 -19950
rect 8300 -20200 11850 -20050
rect 12500 -20050 12550 -19950
rect 13000 -20050 13050 -19950
rect 13500 -20050 13550 -19950
rect 14000 -20050 14050 -19950
rect 14500 -20050 14550 -19950
rect 15000 -20050 15050 -19950
rect 15500 -20050 15550 -19950
rect 16000 -20050 16050 -19950
rect 16500 -20050 16550 -19950
rect 17000 -20050 17050 -19950
rect 17500 -20050 17550 -19950
rect 18000 -20050 18050 -19950
rect 18500 -20050 18550 -19950
rect 19000 -20050 19050 -19950
rect 19500 -20050 19550 -19950
rect 20000 -20050 20050 -19950
rect 12500 -20200 20050 -20050
rect 20700 -20050 20750 -19950
rect 21200 -20050 21250 -19950
rect 21700 -20050 21750 -19950
rect 22200 -20050 22250 -19950
rect 22700 -20050 22750 -19950
rect 23200 -20050 23250 -19950
rect 23700 -20050 23750 -19950
rect 24200 -20050 24250 -19950
rect 20700 -20200 24250 -20050
rect 24900 -20050 24950 -19950
rect 25400 -20050 25450 -19950
rect 25900 -20050 25950 -19950
rect 26400 -20050 26450 -19950
rect 24900 -20200 26450 -20050
rect 27100 -20050 27150 -19950
rect 27600 -20050 27650 -19950
rect 27100 -20200 27650 -20050
rect 28300 -20200 28350 -19950
rect 29000 -20050 29050 -19950
rect 29500 -20050 29550 -19950
rect 30000 -20050 30050 -19950
rect 30500 -20050 30550 -19950
rect 29000 -20200 30550 -20050
rect 31200 -20050 31250 -19950
rect 31700 -20050 31750 -19950
rect 31200 -20200 31750 -20050
rect 32400 -20200 32450 -19950
use cap1  cap1_0
timestamp 1666367459
transform 1 0 36400 0 1 0
box 0 0 350 2250
use cap1  cap1_1
timestamp 1666367459
transform 1 0 40500 0 -1 -995
box 0 0 350 2250
use cap1  cap1_2
timestamp 1666367459
transform 1 0 41200 0 -1 -995
box 0 0 350 2250
use cap1  cap1_3
timestamp 1666367459
transform 1 0 36400 0 -1 -995
box 0 0 350 2250
use cap1  cap1_4
timestamp 1666367459
transform 1 0 41200 0 1 0
box 0 0 350 2250
use cap1  cap1_5
timestamp 1666367459
transform 1 0 40500 0 1 0
box 0 0 350 2250
use cap2  cap2_0
timestamp 1666367418
transform 1 0 35200 0 1 0
box 0 0 850 2250
use cap2  cap2_1
timestamp 1666367418
transform 1 0 39300 0 -1 -995
box 0 0 850 2250
use cap2  cap2_2
timestamp 1666367418
transform 1 0 35200 0 -1 -995
box 0 0 850 2250
use cap2  cap2_3
timestamp 1666367418
transform 1 0 39300 0 1 0
box 0 0 850 2250
use cap4  cap4_0
timestamp 1666367387
transform 1 0 33000 0 1 0
box 0 0 1850 2250
use cap4  cap4_1
timestamp 1666367387
transform 1 0 37100 0 1 0
box 0 0 1850 2250
use cap4  cap4_2
timestamp 1666367387
transform 1 0 37100 0 -1 -995
box 0 0 1850 2250
use cap4  cap4_3
timestamp 1666367387
transform 1 0 33000 0 -1 -995
box 0 0 1850 2250
use cap8  cap8_0
timestamp 1666311562
transform 1 0 28200 0 1 0
box 0 0 350 19005
use cap8  cap8_1
timestamp 1666311562
transform 1 0 32300 0 1 0
box 0 0 350 19005
use cap8  cap8_2
timestamp 1666311562
transform 1 0 32300 0 -1 -995
box 0 0 350 19005
use cap8  cap8_3
timestamp 1666311562
transform 1 0 28200 0 -1 -995
box 0 0 350 19005
use cap16  cap16_0
timestamp 1666311401
transform 1 0 27000 0 1 0
box 0 0 850 19005
use cap16  cap16_1
timestamp 1666311401
transform 1 0 31100 0 1 0
box 0 0 850 19005
use cap16  cap16_2
timestamp 1666311401
transform 1 0 31100 0 -1 -995
box 0 0 850 19005
use cap16  cap16_3
timestamp 1666311401
transform 1 0 27000 0 -1 -995
box 0 0 850 19005
use cap32  cap32_0
timestamp 1666311305
transform 1 0 24800 0 1 0
box 0 0 1850 19005
use cap32  cap32_1
timestamp 1666311305
transform 1 0 28900 0 1 0
box 0 0 1850 19005
use cap32  cap32_2
timestamp 1666311305
transform 1 0 28900 0 -1 -995
box 0 0 1850 19005
use cap32  cap32_3
timestamp 1666311305
transform 1 0 24800 0 -1 -995
box 0 0 1850 19005
use cap64  cap64_0
timestamp 1666313508
transform 1 0 20600 0 1 0
box 0 0 3850 19005
use cap64  cap64_1
timestamp 1666313508
transform 1 0 8200 0 1 0
box 0 0 3850 19005
use cap64  cap64_2
timestamp 1666313508
transform 1 0 20600 0 -1 -995
box 0 0 3850 19005
use cap64  cap64_3
timestamp 1666313508
transform 1 0 8200 0 -1 -995
box 0 0 3850 19005
use cap128  cap128_0
timestamp 1666311401
transform 1 0 0 0 1 0
box 0 0 7850 19005
use cap128  cap128_1
timestamp 1666311401
transform 1 0 12400 0 1 0
box 0 0 7850 19005
use cap128  cap128_2
timestamp 1666311401
transform 1 0 12400 0 -1 -995
box 0 0 7850 19005
use cap128  cap128_3
timestamp 1666311401
transform 1 0 0 0 -1 -995
box 0 0 7850 19005
<< labels >>
rlabel metal4 41300 -3395 41350 -3245 1 sw_sp_n9
port 1 n
rlabel metal4 36500 -3395 36550 -3245 1 sw_sp_n8
port 2 n
rlabel metal4 35300 -3395 35850 -3245 1 sw_sp_n7
port 3 n
rlabel metal4 33100 -3395 34650 -3245 1 sw_sp_n6
port 4 n
rlabel metal4 28300 -20200 28350 -19950 1 sw_sp_n5
port 5 n
rlabel metal4 27100 -20200 27650 -20050 1 sw_sp_n4
port 6 n
rlabel metal4 24900 -20200 26450 -20050 1 sw_sp_n3
port 7 n
rlabel metal4 8300 -20200 11850 -20050 1 sw_sp_n2
port 8 n
rlabel metal4 100 -20200 7650 -20050 1 sw_sp_n1
port 9 n
rlabel metal4 300 -200 41550 -50 1 Vin_p
port 10 n
rlabel metal4 300 -950 41550 -800 1 Vin_n
port 11 n
rlabel metal4 41300 2250 41350 2400 1 sw_sp_p9
port 12 n
rlabel metal4 36500 2250 36550 2400 1 sw_sp_p8
port 13 n
rlabel metal4 35300 2250 35850 2400 1 sw_sp_p7
port 14 n
rlabel metal4 33100 2250 34650 2400 1 sw_sp_p6
port 15 n
rlabel metal4 28300 19000 28350 19200 1 sw_sp_p5
port 16 n
rlabel metal4 27100 19050 27650 19200 1 sw_sp_p4
port 17 n
rlabel metal4 24900 19050 26450 19200 1 sw_sp_p3
port 18 n
rlabel metal4 8300 19050 11850 19200 1 sw_sp_p2
port 19 n
rlabel metal4 100 19050 7650 19200 1 sw_sp_p1
port 20 n
rlabel metal4 40600 2250 40650 2400 1 sw_p8
port 21 n
rlabel metal4 39400 2250 39950 2400 1 sw_p7
port 22 n
rlabel metal4 37200 2250 38750 2400 1 sw_p6
port 23 n
rlabel metal4 32400 19000 32450 19200 1 sw_p5
port 24 n
rlabel metal4 31200 19050 31750 19200 1 sw_p4
port 25 n
rlabel metal4 29000 19050 30550 19200 1 sw_p3
port 26 n
rlabel metal4 20700 19050 24250 19200 1 sw_p2
port 27 n
rlabel metal4 12500 19050 20050 19200 1 sw_p1
port 28 n
rlabel metal4 40600 -3395 40650 -3245 1 sw_n8
port 29 n
rlabel metal4 39400 -3395 39950 -3245 1 sw_n7
port 30 n
rlabel metal4 37200 -3395 38750 -3245 1 sw_n6
port 31 n
rlabel metal4 32400 -20200 32450 -19950 1 sw_n5
port 32 n
rlabel metal4 31200 -20200 31750 -20050 1 sw_n4
port 33 n
rlabel metal4 29000 -20200 30550 -20050 1 sw_n3
port 34 n
rlabel metal4 20700 -20200 24250 -20050 1 sw_n2
port 35 n
rlabel metal4 12500 -20200 20050 -20050 1 sw_n1
port 36 n
<< end >>
