magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -1904 17972 -1132 18000
rect -1904 13738 -1216 17972
rect -1152 13738 -1132 17972
rect -1904 13710 -1132 13738
rect -892 17972 -120 18000
rect -892 13738 -204 17972
rect -140 13738 -120 17972
rect -892 13710 -120 13738
rect 120 17972 892 18000
rect 120 13738 808 17972
rect 872 13738 892 17972
rect 120 13710 892 13738
rect 1132 17972 1904 18000
rect 1132 13738 1820 17972
rect 1884 13738 1904 17972
rect 1132 13710 1904 13738
rect -1904 13442 -1132 13470
rect -1904 9208 -1216 13442
rect -1152 9208 -1132 13442
rect -1904 9180 -1132 9208
rect -892 13442 -120 13470
rect -892 9208 -204 13442
rect -140 9208 -120 13442
rect -892 9180 -120 9208
rect 120 13442 892 13470
rect 120 9208 808 13442
rect 872 9208 892 13442
rect 120 9180 892 9208
rect 1132 13442 1904 13470
rect 1132 9208 1820 13442
rect 1884 9208 1904 13442
rect 1132 9180 1904 9208
rect -1904 8912 -1132 8940
rect -1904 4678 -1216 8912
rect -1152 4678 -1132 8912
rect -1904 4650 -1132 4678
rect -892 8912 -120 8940
rect -892 4678 -204 8912
rect -140 4678 -120 8912
rect -892 4650 -120 4678
rect 120 8912 892 8940
rect 120 4678 808 8912
rect 872 4678 892 8912
rect 120 4650 892 4678
rect 1132 8912 1904 8940
rect 1132 4678 1820 8912
rect 1884 4678 1904 8912
rect 1132 4650 1904 4678
rect -1904 4382 -1132 4410
rect -1904 148 -1216 4382
rect -1152 148 -1132 4382
rect -1904 120 -1132 148
rect -892 4382 -120 4410
rect -892 148 -204 4382
rect -140 148 -120 4382
rect -892 120 -120 148
rect 120 4382 892 4410
rect 120 148 808 4382
rect 872 148 892 4382
rect 120 120 892 148
rect 1132 4382 1904 4410
rect 1132 148 1820 4382
rect 1884 148 1904 4382
rect 1132 120 1904 148
rect -1904 -148 -1132 -120
rect -1904 -4382 -1216 -148
rect -1152 -4382 -1132 -148
rect -1904 -4410 -1132 -4382
rect -892 -148 -120 -120
rect -892 -4382 -204 -148
rect -140 -4382 -120 -148
rect -892 -4410 -120 -4382
rect 120 -148 892 -120
rect 120 -4382 808 -148
rect 872 -4382 892 -148
rect 120 -4410 892 -4382
rect 1132 -148 1904 -120
rect 1132 -4382 1820 -148
rect 1884 -4382 1904 -148
rect 1132 -4410 1904 -4382
rect -1904 -4678 -1132 -4650
rect -1904 -8912 -1216 -4678
rect -1152 -8912 -1132 -4678
rect -1904 -8940 -1132 -8912
rect -892 -4678 -120 -4650
rect -892 -8912 -204 -4678
rect -140 -8912 -120 -4678
rect -892 -8940 -120 -8912
rect 120 -4678 892 -4650
rect 120 -8912 808 -4678
rect 872 -8912 892 -4678
rect 120 -8940 892 -8912
rect 1132 -4678 1904 -4650
rect 1132 -8912 1820 -4678
rect 1884 -8912 1904 -4678
rect 1132 -8940 1904 -8912
rect -1904 -9208 -1132 -9180
rect -1904 -13442 -1216 -9208
rect -1152 -13442 -1132 -9208
rect -1904 -13470 -1132 -13442
rect -892 -9208 -120 -9180
rect -892 -13442 -204 -9208
rect -140 -13442 -120 -9208
rect -892 -13470 -120 -13442
rect 120 -9208 892 -9180
rect 120 -13442 808 -9208
rect 872 -13442 892 -9208
rect 120 -13470 892 -13442
rect 1132 -9208 1904 -9180
rect 1132 -13442 1820 -9208
rect 1884 -13442 1904 -9208
rect 1132 -13470 1904 -13442
rect -1904 -13738 -1132 -13710
rect -1904 -17972 -1216 -13738
rect -1152 -17972 -1132 -13738
rect -1904 -18000 -1132 -17972
rect -892 -13738 -120 -13710
rect -892 -17972 -204 -13738
rect -140 -17972 -120 -13738
rect -892 -18000 -120 -17972
rect 120 -13738 892 -13710
rect 120 -17972 808 -13738
rect 872 -17972 892 -13738
rect 120 -18000 892 -17972
rect 1132 -13738 1904 -13710
rect 1132 -17972 1820 -13738
rect 1884 -17972 1904 -13738
rect 1132 -18000 1904 -17972
<< via3 >>
rect -1216 13738 -1152 17972
rect -204 13738 -140 17972
rect 808 13738 872 17972
rect 1820 13738 1884 17972
rect -1216 9208 -1152 13442
rect -204 9208 -140 13442
rect 808 9208 872 13442
rect 1820 9208 1884 13442
rect -1216 4678 -1152 8912
rect -204 4678 -140 8912
rect 808 4678 872 8912
rect 1820 4678 1884 8912
rect -1216 148 -1152 4382
rect -204 148 -140 4382
rect 808 148 872 4382
rect 1820 148 1884 4382
rect -1216 -4382 -1152 -148
rect -204 -4382 -140 -148
rect 808 -4382 872 -148
rect 1820 -4382 1884 -148
rect -1216 -8912 -1152 -4678
rect -204 -8912 -140 -4678
rect 808 -8912 872 -4678
rect 1820 -8912 1884 -4678
rect -1216 -13442 -1152 -9208
rect -204 -13442 -140 -9208
rect 808 -13442 872 -9208
rect 1820 -13442 1884 -9208
rect -1216 -17972 -1152 -13738
rect -204 -17972 -140 -13738
rect 808 -17972 872 -13738
rect 1820 -17972 1884 -13738
<< mimcap >>
rect -1864 17920 -1464 17960
rect -1864 13790 -1824 17920
rect -1504 13790 -1464 17920
rect -1864 13750 -1464 13790
rect -852 17920 -452 17960
rect -852 13790 -812 17920
rect -492 13790 -452 17920
rect -852 13750 -452 13790
rect 160 17920 560 17960
rect 160 13790 200 17920
rect 520 13790 560 17920
rect 160 13750 560 13790
rect 1172 17920 1572 17960
rect 1172 13790 1212 17920
rect 1532 13790 1572 17920
rect 1172 13750 1572 13790
rect -1864 13390 -1464 13430
rect -1864 9260 -1824 13390
rect -1504 9260 -1464 13390
rect -1864 9220 -1464 9260
rect -852 13390 -452 13430
rect -852 9260 -812 13390
rect -492 9260 -452 13390
rect -852 9220 -452 9260
rect 160 13390 560 13430
rect 160 9260 200 13390
rect 520 9260 560 13390
rect 160 9220 560 9260
rect 1172 13390 1572 13430
rect 1172 9260 1212 13390
rect 1532 9260 1572 13390
rect 1172 9220 1572 9260
rect -1864 8860 -1464 8900
rect -1864 4730 -1824 8860
rect -1504 4730 -1464 8860
rect -1864 4690 -1464 4730
rect -852 8860 -452 8900
rect -852 4730 -812 8860
rect -492 4730 -452 8860
rect -852 4690 -452 4730
rect 160 8860 560 8900
rect 160 4730 200 8860
rect 520 4730 560 8860
rect 160 4690 560 4730
rect 1172 8860 1572 8900
rect 1172 4730 1212 8860
rect 1532 4730 1572 8860
rect 1172 4690 1572 4730
rect -1864 4330 -1464 4370
rect -1864 200 -1824 4330
rect -1504 200 -1464 4330
rect -1864 160 -1464 200
rect -852 4330 -452 4370
rect -852 200 -812 4330
rect -492 200 -452 4330
rect -852 160 -452 200
rect 160 4330 560 4370
rect 160 200 200 4330
rect 520 200 560 4330
rect 160 160 560 200
rect 1172 4330 1572 4370
rect 1172 200 1212 4330
rect 1532 200 1572 4330
rect 1172 160 1572 200
rect -1864 -200 -1464 -160
rect -1864 -4330 -1824 -200
rect -1504 -4330 -1464 -200
rect -1864 -4370 -1464 -4330
rect -852 -200 -452 -160
rect -852 -4330 -812 -200
rect -492 -4330 -452 -200
rect -852 -4370 -452 -4330
rect 160 -200 560 -160
rect 160 -4330 200 -200
rect 520 -4330 560 -200
rect 160 -4370 560 -4330
rect 1172 -200 1572 -160
rect 1172 -4330 1212 -200
rect 1532 -4330 1572 -200
rect 1172 -4370 1572 -4330
rect -1864 -4730 -1464 -4690
rect -1864 -8860 -1824 -4730
rect -1504 -8860 -1464 -4730
rect -1864 -8900 -1464 -8860
rect -852 -4730 -452 -4690
rect -852 -8860 -812 -4730
rect -492 -8860 -452 -4730
rect -852 -8900 -452 -8860
rect 160 -4730 560 -4690
rect 160 -8860 200 -4730
rect 520 -8860 560 -4730
rect 160 -8900 560 -8860
rect 1172 -4730 1572 -4690
rect 1172 -8860 1212 -4730
rect 1532 -8860 1572 -4730
rect 1172 -8900 1572 -8860
rect -1864 -9260 -1464 -9220
rect -1864 -13390 -1824 -9260
rect -1504 -13390 -1464 -9260
rect -1864 -13430 -1464 -13390
rect -852 -9260 -452 -9220
rect -852 -13390 -812 -9260
rect -492 -13390 -452 -9260
rect -852 -13430 -452 -13390
rect 160 -9260 560 -9220
rect 160 -13390 200 -9260
rect 520 -13390 560 -9260
rect 160 -13430 560 -13390
rect 1172 -9260 1572 -9220
rect 1172 -13390 1212 -9260
rect 1532 -13390 1572 -9260
rect 1172 -13430 1572 -13390
rect -1864 -13790 -1464 -13750
rect -1864 -17920 -1824 -13790
rect -1504 -17920 -1464 -13790
rect -1864 -17960 -1464 -17920
rect -852 -13790 -452 -13750
rect -852 -17920 -812 -13790
rect -492 -17920 -452 -13790
rect -852 -17960 -452 -17920
rect 160 -13790 560 -13750
rect 160 -17920 200 -13790
rect 520 -17920 560 -13790
rect 160 -17960 560 -17920
rect 1172 -13790 1572 -13750
rect 1172 -17920 1212 -13790
rect 1532 -17920 1572 -13790
rect 1172 -17960 1572 -17920
<< mimcapcontact >>
rect -1824 13790 -1504 17920
rect -812 13790 -492 17920
rect 200 13790 520 17920
rect 1212 13790 1532 17920
rect -1824 9260 -1504 13390
rect -812 9260 -492 13390
rect 200 9260 520 13390
rect 1212 9260 1532 13390
rect -1824 4730 -1504 8860
rect -812 4730 -492 8860
rect 200 4730 520 8860
rect 1212 4730 1532 8860
rect -1824 200 -1504 4330
rect -812 200 -492 4330
rect 200 200 520 4330
rect 1212 200 1532 4330
rect -1824 -4330 -1504 -200
rect -812 -4330 -492 -200
rect 200 -4330 520 -200
rect 1212 -4330 1532 -200
rect -1824 -8860 -1504 -4730
rect -812 -8860 -492 -4730
rect 200 -8860 520 -4730
rect 1212 -8860 1532 -4730
rect -1824 -13390 -1504 -9260
rect -812 -13390 -492 -9260
rect 200 -13390 520 -9260
rect 1212 -13390 1532 -9260
rect -1824 -17920 -1504 -13790
rect -812 -17920 -492 -13790
rect 200 -17920 520 -13790
rect 1212 -17920 1532 -13790
<< metal4 >>
rect -1716 17921 -1612 18120
rect -1236 17972 -1132 18120
rect -1825 17920 -1503 17921
rect -1825 13790 -1824 17920
rect -1504 13790 -1503 17920
rect -1825 13789 -1503 13790
rect -1716 13391 -1612 13789
rect -1236 13738 -1216 17972
rect -1152 13738 -1132 17972
rect -704 17921 -600 18120
rect -224 17972 -120 18120
rect -813 17920 -491 17921
rect -813 13790 -812 17920
rect -492 13790 -491 17920
rect -813 13789 -491 13790
rect -1236 13442 -1132 13738
rect -1825 13390 -1503 13391
rect -1825 9260 -1824 13390
rect -1504 9260 -1503 13390
rect -1825 9259 -1503 9260
rect -1716 8861 -1612 9259
rect -1236 9208 -1216 13442
rect -1152 9208 -1132 13442
rect -704 13391 -600 13789
rect -224 13738 -204 17972
rect -140 13738 -120 17972
rect 308 17921 412 18120
rect 788 17972 892 18120
rect 199 17920 521 17921
rect 199 13790 200 17920
rect 520 13790 521 17920
rect 199 13789 521 13790
rect -224 13442 -120 13738
rect -813 13390 -491 13391
rect -813 9260 -812 13390
rect -492 9260 -491 13390
rect -813 9259 -491 9260
rect -1236 8912 -1132 9208
rect -1825 8860 -1503 8861
rect -1825 4730 -1824 8860
rect -1504 4730 -1503 8860
rect -1825 4729 -1503 4730
rect -1716 4331 -1612 4729
rect -1236 4678 -1216 8912
rect -1152 4678 -1132 8912
rect -704 8861 -600 9259
rect -224 9208 -204 13442
rect -140 9208 -120 13442
rect 308 13391 412 13789
rect 788 13738 808 17972
rect 872 13738 892 17972
rect 1320 17921 1424 18120
rect 1800 17972 1904 18120
rect 1211 17920 1533 17921
rect 1211 13790 1212 17920
rect 1532 13790 1533 17920
rect 1211 13789 1533 13790
rect 788 13442 892 13738
rect 199 13390 521 13391
rect 199 9260 200 13390
rect 520 9260 521 13390
rect 199 9259 521 9260
rect -224 8912 -120 9208
rect -813 8860 -491 8861
rect -813 4730 -812 8860
rect -492 4730 -491 8860
rect -813 4729 -491 4730
rect -1236 4382 -1132 4678
rect -1825 4330 -1503 4331
rect -1825 200 -1824 4330
rect -1504 200 -1503 4330
rect -1825 199 -1503 200
rect -1716 -199 -1612 199
rect -1236 148 -1216 4382
rect -1152 148 -1132 4382
rect -704 4331 -600 4729
rect -224 4678 -204 8912
rect -140 4678 -120 8912
rect 308 8861 412 9259
rect 788 9208 808 13442
rect 872 9208 892 13442
rect 1320 13391 1424 13789
rect 1800 13738 1820 17972
rect 1884 13738 1904 17972
rect 1800 13442 1904 13738
rect 1211 13390 1533 13391
rect 1211 9260 1212 13390
rect 1532 9260 1533 13390
rect 1211 9259 1533 9260
rect 788 8912 892 9208
rect 199 8860 521 8861
rect 199 4730 200 8860
rect 520 4730 521 8860
rect 199 4729 521 4730
rect -224 4382 -120 4678
rect -813 4330 -491 4331
rect -813 200 -812 4330
rect -492 200 -491 4330
rect -813 199 -491 200
rect -1236 -148 -1132 148
rect -1825 -200 -1503 -199
rect -1825 -4330 -1824 -200
rect -1504 -4330 -1503 -200
rect -1825 -4331 -1503 -4330
rect -1716 -4729 -1612 -4331
rect -1236 -4382 -1216 -148
rect -1152 -4382 -1132 -148
rect -704 -199 -600 199
rect -224 148 -204 4382
rect -140 148 -120 4382
rect 308 4331 412 4729
rect 788 4678 808 8912
rect 872 4678 892 8912
rect 1320 8861 1424 9259
rect 1800 9208 1820 13442
rect 1884 9208 1904 13442
rect 1800 8912 1904 9208
rect 1211 8860 1533 8861
rect 1211 4730 1212 8860
rect 1532 4730 1533 8860
rect 1211 4729 1533 4730
rect 788 4382 892 4678
rect 199 4330 521 4331
rect 199 200 200 4330
rect 520 200 521 4330
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -4330 -812 -200
rect -492 -4330 -491 -200
rect -813 -4331 -491 -4330
rect -1236 -4678 -1132 -4382
rect -1825 -4730 -1503 -4729
rect -1825 -8860 -1824 -4730
rect -1504 -8860 -1503 -4730
rect -1825 -8861 -1503 -8860
rect -1716 -9259 -1612 -8861
rect -1236 -8912 -1216 -4678
rect -1152 -8912 -1132 -4678
rect -704 -4729 -600 -4331
rect -224 -4382 -204 -148
rect -140 -4382 -120 -148
rect 308 -199 412 199
rect 788 148 808 4382
rect 872 148 892 4382
rect 1320 4331 1424 4729
rect 1800 4678 1820 8912
rect 1884 4678 1904 8912
rect 1800 4382 1904 4678
rect 1211 4330 1533 4331
rect 1211 200 1212 4330
rect 1532 200 1533 4330
rect 1211 199 1533 200
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -4330 200 -200
rect 520 -4330 521 -200
rect 199 -4331 521 -4330
rect -224 -4678 -120 -4382
rect -813 -4730 -491 -4729
rect -813 -8860 -812 -4730
rect -492 -8860 -491 -4730
rect -813 -8861 -491 -8860
rect -1236 -9208 -1132 -8912
rect -1825 -9260 -1503 -9259
rect -1825 -13390 -1824 -9260
rect -1504 -13390 -1503 -9260
rect -1825 -13391 -1503 -13390
rect -1716 -13789 -1612 -13391
rect -1236 -13442 -1216 -9208
rect -1152 -13442 -1132 -9208
rect -704 -9259 -600 -8861
rect -224 -8912 -204 -4678
rect -140 -8912 -120 -4678
rect 308 -4729 412 -4331
rect 788 -4382 808 -148
rect 872 -4382 892 -148
rect 1320 -199 1424 199
rect 1800 148 1820 4382
rect 1884 148 1904 4382
rect 1800 -148 1904 148
rect 1211 -200 1533 -199
rect 1211 -4330 1212 -200
rect 1532 -4330 1533 -200
rect 1211 -4331 1533 -4330
rect 788 -4678 892 -4382
rect 199 -4730 521 -4729
rect 199 -8860 200 -4730
rect 520 -8860 521 -4730
rect 199 -8861 521 -8860
rect -224 -9208 -120 -8912
rect -813 -9260 -491 -9259
rect -813 -13390 -812 -9260
rect -492 -13390 -491 -9260
rect -813 -13391 -491 -13390
rect -1236 -13738 -1132 -13442
rect -1825 -13790 -1503 -13789
rect -1825 -17920 -1824 -13790
rect -1504 -17920 -1503 -13790
rect -1825 -17921 -1503 -17920
rect -1716 -18120 -1612 -17921
rect -1236 -17972 -1216 -13738
rect -1152 -17972 -1132 -13738
rect -704 -13789 -600 -13391
rect -224 -13442 -204 -9208
rect -140 -13442 -120 -9208
rect 308 -9259 412 -8861
rect 788 -8912 808 -4678
rect 872 -8912 892 -4678
rect 1320 -4729 1424 -4331
rect 1800 -4382 1820 -148
rect 1884 -4382 1904 -148
rect 1800 -4678 1904 -4382
rect 1211 -4730 1533 -4729
rect 1211 -8860 1212 -4730
rect 1532 -8860 1533 -4730
rect 1211 -8861 1533 -8860
rect 788 -9208 892 -8912
rect 199 -9260 521 -9259
rect 199 -13390 200 -9260
rect 520 -13390 521 -9260
rect 199 -13391 521 -13390
rect -224 -13738 -120 -13442
rect -813 -13790 -491 -13789
rect -813 -17920 -812 -13790
rect -492 -17920 -491 -13790
rect -813 -17921 -491 -17920
rect -1236 -18120 -1132 -17972
rect -704 -18120 -600 -17921
rect -224 -17972 -204 -13738
rect -140 -17972 -120 -13738
rect 308 -13789 412 -13391
rect 788 -13442 808 -9208
rect 872 -13442 892 -9208
rect 1320 -9259 1424 -8861
rect 1800 -8912 1820 -4678
rect 1884 -8912 1904 -4678
rect 1800 -9208 1904 -8912
rect 1211 -9260 1533 -9259
rect 1211 -13390 1212 -9260
rect 1532 -13390 1533 -9260
rect 1211 -13391 1533 -13390
rect 788 -13738 892 -13442
rect 199 -13790 521 -13789
rect 199 -17920 200 -13790
rect 520 -17920 521 -13790
rect 199 -17921 521 -17920
rect -224 -18120 -120 -17972
rect 308 -18120 412 -17921
rect 788 -17972 808 -13738
rect 872 -17972 892 -13738
rect 1320 -13789 1424 -13391
rect 1800 -13442 1820 -9208
rect 1884 -13442 1904 -9208
rect 1800 -13738 1904 -13442
rect 1211 -13790 1533 -13789
rect 1211 -17920 1212 -13790
rect 1532 -17920 1533 -13790
rect 1211 -17921 1533 -17920
rect 788 -18120 892 -17972
rect 1320 -18120 1424 -17921
rect 1800 -17972 1820 -13738
rect 1884 -17972 1904 -13738
rect 1800 -18120 1904 -17972
<< properties >>
string FIXED_BBOX 1132 13710 1612 18000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
