magic
tech sky130A
magscale 1 2
timestamp 1666807393
<< error_p >>
rect -269 163 -211 169
rect -77 163 -19 169
rect 115 163 173 169
rect 307 163 365 169
rect -269 129 -257 163
rect -77 129 -65 163
rect 115 129 127 163
rect 307 129 319 163
rect -269 123 -211 129
rect -77 123 -19 129
rect 115 123 173 129
rect 307 123 365 129
rect -365 -129 -307 -123
rect -173 -129 -115 -123
rect 19 -129 77 -123
rect 211 -129 269 -123
rect -365 -163 -353 -129
rect -173 -163 -161 -129
rect 19 -163 31 -129
rect 211 -163 223 -129
rect -365 -169 -307 -163
rect -173 -169 -115 -163
rect 19 -169 77 -163
rect 211 -169 269 -163
<< nmos >>
rect -351 -91 -321 91
rect -255 -91 -225 91
rect -159 -91 -129 91
rect -63 -91 -33 91
rect 33 -91 63 91
rect 129 -91 159 91
rect 225 -91 255 91
rect 321 -91 351 91
<< ndiff >>
rect -413 79 -351 91
rect -413 -79 -401 79
rect -367 -79 -351 79
rect -413 -91 -351 -79
rect -321 79 -255 91
rect -321 -79 -305 79
rect -271 -79 -255 79
rect -321 -91 -255 -79
rect -225 79 -159 91
rect -225 -79 -209 79
rect -175 -79 -159 79
rect -225 -91 -159 -79
rect -129 79 -63 91
rect -129 -79 -113 79
rect -79 -79 -63 79
rect -129 -91 -63 -79
rect -33 79 33 91
rect -33 -79 -17 79
rect 17 -79 33 79
rect -33 -91 33 -79
rect 63 79 129 91
rect 63 -79 79 79
rect 113 -79 129 79
rect 63 -91 129 -79
rect 159 79 225 91
rect 159 -79 175 79
rect 209 -79 225 79
rect 159 -91 225 -79
rect 255 79 321 91
rect 255 -79 271 79
rect 305 -79 321 79
rect 255 -91 321 -79
rect 351 79 413 91
rect 351 -79 367 79
rect 401 -79 413 79
rect 351 -91 413 -79
<< ndiffc >>
rect -401 -79 -367 79
rect -305 -79 -271 79
rect -209 -79 -175 79
rect -113 -79 -79 79
rect -17 -79 17 79
rect 79 -79 113 79
rect 175 -79 209 79
rect 271 -79 305 79
rect 367 -79 401 79
<< poly >>
rect -273 163 -207 179
rect -273 129 -257 163
rect -223 129 -207 163
rect -351 91 -321 117
rect -273 113 -207 129
rect -81 163 -15 179
rect -81 129 -65 163
rect -31 129 -15 163
rect -255 91 -225 113
rect -159 91 -129 117
rect -81 113 -15 129
rect 111 163 177 179
rect 111 129 127 163
rect 161 129 177 163
rect -63 91 -33 113
rect 33 91 63 117
rect 111 113 177 129
rect 303 163 369 179
rect 303 129 319 163
rect 353 129 369 163
rect 129 91 159 113
rect 225 91 255 117
rect 303 113 369 129
rect 321 91 351 113
rect -351 -113 -321 -91
rect -369 -129 -303 -113
rect -255 -117 -225 -91
rect -159 -113 -129 -91
rect -369 -163 -353 -129
rect -319 -163 -303 -129
rect -369 -179 -303 -163
rect -177 -129 -111 -113
rect -63 -117 -33 -91
rect 33 -113 63 -91
rect -177 -163 -161 -129
rect -127 -163 -111 -129
rect -177 -179 -111 -163
rect 15 -129 81 -113
rect 129 -117 159 -91
rect 225 -113 255 -91
rect 15 -163 31 -129
rect 65 -163 81 -129
rect 15 -179 81 -163
rect 207 -129 273 -113
rect 321 -117 351 -91
rect 207 -163 223 -129
rect 257 -163 273 -129
rect 207 -179 273 -163
<< polycont >>
rect -257 129 -223 163
rect -65 129 -31 163
rect 127 129 161 163
rect 319 129 353 163
rect -353 -163 -319 -129
rect -161 -163 -127 -129
rect 31 -163 65 -129
rect 223 -163 257 -129
<< locali >>
rect -273 129 -257 163
rect -223 129 -207 163
rect -81 129 -65 163
rect -31 129 -15 163
rect 111 129 127 163
rect 161 129 177 163
rect 303 129 319 163
rect 353 129 369 163
rect -401 79 -367 95
rect -401 -95 -367 -79
rect -305 79 -271 95
rect -305 -95 -271 -79
rect -209 79 -175 95
rect -209 -95 -175 -79
rect -113 79 -79 95
rect -113 -95 -79 -79
rect -17 79 17 95
rect -17 -95 17 -79
rect 79 79 113 95
rect 79 -95 113 -79
rect 175 79 209 95
rect 175 -95 209 -79
rect 271 79 305 95
rect 271 -95 305 -79
rect 367 79 401 95
rect 367 -95 401 -79
rect -369 -163 -353 -129
rect -319 -163 -303 -129
rect -177 -163 -161 -129
rect -127 -163 -111 -129
rect 15 -163 31 -129
rect 65 -163 81 -129
rect 207 -163 223 -129
rect 257 -163 273 -129
<< viali >>
rect -257 129 -223 163
rect -65 129 -31 163
rect 127 129 161 163
rect 319 129 353 163
rect -401 -79 -367 79
rect -305 -62 -271 -7
rect -209 -79 -175 79
rect -113 -62 -79 -7
rect -17 -79 17 79
rect 79 -62 113 -7
rect 175 -79 209 79
rect 271 -62 305 -7
rect 367 -79 401 79
rect -353 -163 -319 -129
rect -161 -163 -127 -129
rect 31 -163 65 -129
rect 223 -163 257 -129
<< metal1 >>
rect -269 163 -211 169
rect -269 129 -257 163
rect -223 129 -211 163
rect -269 123 -211 129
rect -77 163 -19 169
rect -77 129 -65 163
rect -31 129 -19 163
rect -77 123 -19 129
rect 115 163 173 169
rect 115 129 127 163
rect 161 129 173 163
rect 115 123 173 129
rect 307 163 365 169
rect 307 129 319 163
rect 353 129 365 163
rect 307 123 365 129
rect -407 79 -361 91
rect -407 -79 -401 79
rect -367 -79 -361 79
rect -215 79 -169 91
rect -311 -7 -265 5
rect -311 -62 -305 -7
rect -271 -62 -265 -7
rect -311 -74 -265 -62
rect -407 -91 -361 -79
rect -215 -79 -209 79
rect -175 -79 -169 79
rect -23 79 23 91
rect -119 -7 -73 5
rect -119 -62 -113 -7
rect -79 -62 -73 -7
rect -119 -74 -73 -62
rect -215 -91 -169 -79
rect -23 -79 -17 79
rect 17 -79 23 79
rect 169 79 215 91
rect 73 -7 119 5
rect 73 -62 79 -7
rect 113 -62 119 -7
rect 73 -74 119 -62
rect -23 -91 23 -79
rect 169 -79 175 79
rect 209 -79 215 79
rect 361 79 407 91
rect 265 -7 311 5
rect 265 -62 271 -7
rect 305 -62 311 -7
rect 265 -74 311 -62
rect 169 -91 215 -79
rect 361 -79 367 79
rect 401 -79 407 79
rect 361 -91 407 -79
rect -365 -129 -307 -123
rect -365 -163 -353 -129
rect -319 -163 -307 -129
rect -365 -169 -307 -163
rect -173 -129 -115 -123
rect -173 -163 -161 -129
rect -127 -163 -115 -129
rect -173 -169 -115 -163
rect 19 -129 77 -123
rect 19 -163 31 -129
rect 65 -163 77 -129
rect 19 -169 77 -163
rect 211 -129 269 -123
rect 211 -163 223 -129
rect 257 -163 269 -129
rect 211 -169 269 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +35 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
