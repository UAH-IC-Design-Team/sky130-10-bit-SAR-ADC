magic
tech sky130A
magscale 1 2
timestamp 1667500811
<< error_s >>
rect 10998 7400 11740 7574
rect 12000 7400 12734 7574
rect 11990 6954 11996 7320
rect 11252 6800 11742 6954
rect 11990 6800 12480 6954
rect 9610 6758 9656 6770
rect 14120 6758 14166 6770
rect 9610 6724 9616 6758
rect 14120 6724 14126 6758
rect 9610 6712 9656 6724
rect 14120 6712 14166 6724
rect 10720 6662 10766 6674
rect 13010 6662 13056 6674
rect 10720 6628 10726 6662
rect 13010 6628 13016 6662
rect 10720 6616 10766 6628
rect 13010 6616 13056 6628
rect 9610 6566 9656 6578
rect 14120 6566 14166 6578
rect 9610 6532 9616 6566
rect 14120 6532 14126 6566
rect 9610 6520 9656 6532
rect 14120 6520 14166 6532
rect 10720 6470 10766 6482
rect 13010 6470 13056 6482
rect 10720 6436 10726 6470
rect 13010 6436 13016 6470
rect 10720 6424 10766 6436
rect 13010 6424 13056 6436
rect 9610 6374 9656 6386
rect 14120 6374 14166 6386
rect 9610 6340 9616 6374
rect 14120 6340 14126 6374
rect 9610 6328 9656 6340
rect 14120 6328 14166 6340
rect 10720 6278 10766 6290
rect 13010 6278 13056 6290
rect 10720 6244 10726 6278
rect 13010 6244 13016 6278
rect 10720 6232 10766 6244
rect 13010 6232 13056 6244
rect 9610 6182 9656 6194
rect 14120 6182 14166 6194
rect 9610 6148 9616 6182
rect 14120 6148 14126 6182
rect 9610 6136 9656 6148
rect 14120 6136 14166 6148
rect 10720 6086 10766 6098
rect 13010 6086 13056 6098
rect 10720 6052 10726 6086
rect 13010 6052 13016 6086
rect 10720 6040 10766 6052
rect 13010 6040 13056 6052
rect 9610 5990 9656 6002
rect 14120 5990 14166 6002
rect 9610 5956 9616 5990
rect 14120 5956 14126 5990
rect 9610 5944 9656 5956
rect 14120 5944 14166 5956
rect 10720 5894 10766 5906
rect 13010 5894 13056 5906
rect 10720 5860 10726 5894
rect 13010 5860 13016 5894
rect 10720 5848 10766 5860
rect 13010 5848 13056 5860
rect 10610 5582 10656 5594
rect 11210 5582 11256 5594
rect 12302 5582 12348 5594
rect 12902 5582 12948 5594
rect 10610 5548 10616 5582
rect 11210 5548 11216 5582
rect 12302 5548 12308 5582
rect 12902 5548 12908 5582
rect 10610 5536 10656 5548
rect 11210 5536 11256 5548
rect 12302 5536 12348 5548
rect 12902 5536 12948 5548
rect 10902 5486 10948 5498
rect 11502 5486 11548 5498
rect 12010 5486 12056 5498
rect 12610 5486 12656 5498
rect 10902 5452 10908 5486
rect 11502 5452 11508 5486
rect 12010 5452 12016 5486
rect 12610 5452 12616 5486
rect 10902 5440 10948 5452
rect 11502 5440 11548 5452
rect 12010 5440 12056 5452
rect 12610 5440 12656 5452
rect 10610 5390 10656 5402
rect 11210 5390 11256 5402
rect 12302 5390 12348 5402
rect 12902 5390 12948 5402
rect 10610 5356 10616 5390
rect 11210 5356 11216 5390
rect 12302 5356 12308 5390
rect 12902 5356 12908 5390
rect 10610 5344 10656 5356
rect 11210 5344 11256 5356
rect 12302 5344 12348 5356
rect 12902 5344 12948 5356
rect 10902 5294 10948 5306
rect 11502 5294 11548 5306
rect 12010 5294 12056 5306
rect 12610 5294 12656 5306
rect 10902 5260 10908 5294
rect 11502 5260 11508 5294
rect 12010 5260 12016 5294
rect 12610 5260 12616 5294
rect 10902 5248 10948 5260
rect 11502 5248 11548 5260
rect 12010 5248 12056 5260
rect 12610 5248 12656 5260
rect 12920 4878 12966 4890
rect 12920 4844 12926 4878
rect 12920 4832 12966 4844
rect 10810 4782 10856 4794
rect 10810 4748 10816 4782
rect 10810 4736 10856 4748
rect 12920 4686 12966 4698
rect 12920 4652 12926 4686
rect 12920 4640 12966 4652
rect 10810 4590 10856 4602
rect 10810 4556 10816 4590
rect 10810 4544 10856 4556
rect 12920 4494 12966 4506
rect 12920 4460 12926 4494
rect 12920 4448 12966 4460
rect 5465 124 5506 130
rect 6055 76 6068 108
rect 7511 -20 7552 -14
rect 8101 -68 8114 -36
rect 9557 -164 9598 -158
rect 10737 -260 10778 -228
rect 12599 -404 12638 -372
rect 13005 -452 13046 -420
rect 13595 -500 13608 -468
use sky130_fd_pr__pfet_01v8_FBQ47L  XM1
timestamp 1666924120
transform 0 1 12600 1 0 7561
box -161 -600 169 560
use sky130_fd_pr__pfet_01v8_5AQ4BN  XM2
timestamp 1666923623
transform 0 -1 11120 1 0 7561
box -161 -620 179 560
use sky130_fd_pr__nfet_01v8_HE67PR  XM3
timestamp 1666918578
transform 0 -1 10188 1 0 6309
box -509 -588 509 588
use sky130_fd_pr__nfet_01v8_HEP4KS  XM4
timestamp 1666918578
transform 0 1 13588 1 0 6309
box -509 -588 509 588
use sky130_fd_pr__nfet_01v8_HZDS97  XM9
timestamp 1666918452
transform 0 -1 11888 1 0 4669
box -269 -1088 269 1088
use sky130_fd_pr__nfet_01v8_9NW33M  XM11
timestamp 1666918578
transform 0 1 12779 1 0 5421
box -221 -179 221 179
use sky130_fd_pr__nfet_01v8_9NW33M  XM12
timestamp 1666918578
transform 0 1 12179 1 0 5421
box -221 -179 221 179
use sky130_fd_pr__nfet_01v8_9NW33M  XM13
timestamp 1666918578
transform 0 -1 11379 1 0 5421
box -221 -179 221 179
use sky130_fd_pr__nfet_01v8_9NW33M  sky130_fd_pr__nfet_01v8_9NW33M_0
timestamp 1666918578
transform 0 -1 10779 1 0 5421
box -221 -179 221 179
use sky130_fd_pr__pfet_01v8_QPTUVJ  sky130_fd_pr__pfet_01v8_QPTUVJ_0
timestamp 1667435677
transform 0 -1 11471 1 0 7057
box -257 -271 263 219
use sky130_fd_pr__pfet_01v8_QPTUVJ  sky130_fd_pr__pfet_01v8_QPTUVJ_1
timestamp 1667435677
transform 0 1 12261 1 0 7057
box -257 -271 263 219
use sky130_fd_pr__pfet_01v8_RPBXXN  sky130_fd_pr__pfet_01v8_RPBXXN_0
timestamp 1666924247
transform 0 -1 12261 -1 0 6249
box -451 -269 449 221
use sky130_fd_pr__pfet_01v8_RPBXXN  sky130_fd_pr__pfet_01v8_RPBXXN_1
timestamp 1666924247
transform 0 1 11461 -1 0 6249
box -451 -269 449 221
use sky130_fd_sc_hd__buf_1  x1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5189 0 1 -89
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5503 0 1 -137
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6093 0 1 -185
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x4
timestamp 1662439860
transform 1 0 7235 0 1 -233
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x5
timestamp 1662439860
transform 1 0 7549 0 1 -281
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x6
timestamp 1662439860
transform 1 0 8139 0 1 -329
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x7
timestamp 1662439860
transform 1 0 9281 0 1 -377
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9595 0 1 -425
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 10369 0 1 -473
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x10
timestamp 1662439860
transform 1 0 10775 0 1 -521
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 11549 0 1 -569
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x12
timestamp 1662439860
transform 1 0 12637 0 1 -665
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  x13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 12323 0 1 -617
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x14
timestamp 1662439860
transform 1 0 13043 0 1 -713
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x15
timestamp 1662439860
transform 1 0 13633 0 1 -761
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  x16
timestamp 1662439860
transform 1 0 14775 0 1 -809
box -38 -48 590 592
<< end >>
