magic
tech sky130A
magscale 1 2
timestamp 1665779562
<< error_p >>
rect -29 626 29 632
rect -29 592 -17 626
rect -29 586 29 592
rect -29 -592 29 -586
rect -29 -626 -17 -592
rect -29 -632 29 -626
<< nwell >>
rect -109 -645 109 645
<< pmos >>
rect -15 -545 15 545
<< pdiff >>
rect -73 533 -15 545
rect -73 -533 -61 533
rect -27 -533 -15 533
rect -73 -545 -15 -533
rect 15 533 73 545
rect 15 -533 27 533
rect 61 -533 73 533
rect 15 -545 73 -533
<< pdiffc >>
rect -61 -533 -27 533
rect 27 -533 61 533
<< poly >>
rect -33 626 33 642
rect -33 592 -17 626
rect 17 592 33 626
rect -33 576 33 592
rect -15 545 15 576
rect -15 -576 15 -545
rect -33 -592 33 -576
rect -33 -626 -17 -592
rect 17 -626 33 -592
rect -33 -642 33 -626
<< polycont >>
rect -17 592 17 626
rect -17 -626 17 -592
<< locali >>
rect -33 592 -17 626
rect 17 592 33 626
rect -61 533 -27 549
rect -61 -549 -27 -533
rect 27 533 61 549
rect 27 -549 61 -533
rect -33 -626 -17 -592
rect 17 -626 33 -592
<< viali >>
rect -17 592 17 626
rect -61 -533 -27 533
rect 27 -533 61 533
rect -17 -626 17 -592
<< metal1 >>
rect -29 626 29 632
rect -29 592 -17 626
rect 17 592 29 626
rect -29 586 29 592
rect -67 533 -21 545
rect -67 -533 -61 533
rect -27 -533 -21 533
rect -67 -545 -21 -533
rect 21 533 67 545
rect 21 -533 27 533
rect 61 -533 67 533
rect 21 -545 67 -533
rect -29 -592 29 -586
rect -29 -626 -17 -592
rect 17 -626 29 -592
rect -29 -632 29 -626
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.445 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
