magic
tech sky130A
magscale 1 2
timestamp 1667690749
<< nwell >>
rect 10520 8460 11520 8800
rect 10660 7540 13070 8080
rect 7730 6100 8510 6110
rect 7730 6080 8620 6100
rect 7731 5834 8620 6080
rect 8841 5900 9780 6110
rect 7730 5779 8620 5834
rect 8840 5779 9780 5900
rect 11060 5800 12680 7280
rect 14180 5780 16410 6110
rect 14190 5779 14442 5780
rect 14550 5779 14796 5780
rect 15190 5779 15432 5780
rect 7320 5080 10240 5410
rect 8110 5079 8356 5080
rect 8930 5079 9176 5080
rect 9750 5079 10398 5080
rect 7540 4370 10150 4710
<< nsubdiff >>
rect 11500 7580 11530 7700
rect 11680 7580 11710 7700
rect 12040 7580 12070 7700
rect 12220 7580 12250 7700
rect 11120 7070 11240 7100
rect 11120 6940 11240 6970
rect 12520 7070 12640 7100
rect 12520 6940 12640 6970
rect 11120 6830 11240 6860
rect 11120 6700 11240 6730
rect 12520 6830 12640 6860
rect 12520 6700 12640 6730
<< nsubdiffcont >>
rect 11530 7580 11680 7700
rect 12070 7580 12220 7700
rect 11120 6970 11240 7070
rect 12520 6970 12640 7070
rect 11120 6730 11240 6830
rect 12520 6730 12640 6830
<< locali >>
rect 10469 8466 10645 8473
rect 10469 8428 10478 8466
rect 10532 8428 10572 8466
rect 10469 8427 10572 8428
rect 10637 8427 10645 8466
rect 10469 8423 10645 8427
rect 10706 8423 10962 8471
rect 11510 7580 11530 7700
rect 11680 7580 11700 7700
rect 12050 7580 12070 7700
rect 12220 7580 12240 7700
rect 11120 7070 11240 7090
rect 11120 6950 11240 6970
rect 12520 7070 12640 7090
rect 12520 6950 12640 6970
rect 11120 6830 11240 6850
rect 11120 6710 11240 6730
rect 12520 6830 12640 6850
rect 12520 6710 12640 6730
rect 8312 5733 8830 5773
rect 9106 5733 9340 5780
rect 14500 5733 14652 5781
rect 15000 5733 15490 5773
rect 8031 5029 8290 5083
rect 8851 5033 9105 5076
rect 9670 5013 9910 5090
rect 9670 5010 9679 5013
rect 7703 4315 7853 4389
rect 9760 4384 9807 4390
rect 8076 4337 8312 4381
rect 8670 4333 9148 4373
rect 9760 4325 9766 4384
rect 9800 4381 9807 4384
rect 9800 4373 9920 4381
rect 9800 4339 9839 4373
rect 9904 4339 9920 4373
rect 9800 4329 9920 4339
rect 9800 4325 9807 4329
rect 9760 4320 9807 4325
<< viali >>
rect 10478 8428 10532 8466
rect 10572 8427 10637 8466
rect 11233 8470 11313 8520
rect 11233 8362 11313 8412
rect 11530 7580 11680 7700
rect 12070 7580 12220 7700
rect 11120 6970 11240 7070
rect 12520 6970 12640 7070
rect 11120 6730 11240 6830
rect 12520 6730 12640 6830
rect 7660 5791 7698 5830
rect 16122 5794 16159 5833
rect 9480 5720 9540 5780
rect 14285 5719 14340 5780
rect 7659 5673 7697 5712
rect 16122 5679 16159 5718
rect 10037 5232 10071 5266
rect 10037 5158 10071 5192
rect 7382 5033 7463 5075
rect 10038 4919 10072 4953
rect 7484 4319 7541 4383
rect 9766 4325 9800 4384
rect 9839 4339 9904 4373
<< metal1 >>
rect 10550 8700 12170 8800
rect 11220 8520 11960 8530
rect 10300 8500 10660 8510
rect 10300 8390 10320 8500
rect 10410 8390 10440 8500
rect 10530 8466 10560 8500
rect 10532 8428 10560 8466
rect 10530 8390 10560 8428
rect 10650 8390 10660 8500
rect 10300 8380 10660 8390
rect 11220 8470 11233 8520
rect 11313 8470 11960 8520
rect 11220 8412 11960 8470
rect 11220 8362 11233 8412
rect 11313 8362 11960 8412
rect 11220 8350 11960 8362
rect 10550 8250 11650 8260
rect 10550 8170 10560 8250
rect 10640 8170 10670 8250
rect 10750 8170 10780 8250
rect 10860 8170 11650 8250
rect 10550 8160 11650 8170
rect 10700 7770 11150 8020
rect 10700 7130 11030 7770
rect 11520 7700 11690 7930
rect 11760 7820 11960 8350
rect 12060 7930 12170 8700
rect 11520 7580 11530 7700
rect 11680 7580 11690 7700
rect 11520 7410 11690 7580
rect 12060 7700 12230 7930
rect 12570 7770 13050 8020
rect 12060 7580 12070 7700
rect 12220 7580 12230 7700
rect 12060 7410 12230 7580
rect 9780 6120 9860 7080
rect 7458 6100 9740 6110
rect 7458 6020 8280 6100
rect 8350 6020 8380 6100
rect 8450 6020 8480 6100
rect 8550 6020 9460 6100
rect 9530 6020 9560 6100
rect 9630 6020 9660 6100
rect 9730 6020 9740 6100
rect 7458 6014 9740 6020
rect 9910 5870 10330 7020
rect 10470 6630 11030 7130
rect 11110 7400 12650 7410
rect 11110 7280 11700 7400
rect 11780 7280 11810 7400
rect 11940 7280 11970 7400
rect 12050 7280 12650 7400
rect 11110 7270 12650 7280
rect 11110 7070 11250 7270
rect 11110 6970 11120 7070
rect 11240 6970 11250 7070
rect 11110 6830 11250 6970
rect 11110 6730 11120 6830
rect 11240 6730 11250 6830
rect 11110 6710 11250 6730
rect 10470 6520 11330 6630
rect 10470 6210 11030 6520
rect 10470 6110 11330 6210
rect 11380 5940 11510 7230
rect 11550 6890 11670 7270
rect 11730 6770 11820 7190
rect 11930 7090 12020 7190
rect 11930 7020 11940 7090
rect 12010 7020 12020 7090
rect 11930 6910 12020 7020
rect 11930 6840 11940 6910
rect 12010 6840 12020 6910
rect 12080 6890 12200 7270
rect 11930 6810 12020 6840
rect 11730 6690 12200 6770
rect 11550 6670 11680 6680
rect 11550 6610 11590 6670
rect 11650 6610 11680 6670
rect 11550 6570 11680 6610
rect 11550 6510 11590 6570
rect 11650 6510 11680 6570
rect 11550 6470 11680 6510
rect 11550 6410 11590 6470
rect 11650 6410 11680 6470
rect 7650 5830 7710 5850
rect 7650 5791 7660 5830
rect 7698 5791 7710 5830
rect 7650 5712 7710 5791
rect 7650 5673 7659 5712
rect 7697 5673 7710 5712
rect 9460 5810 9570 5820
rect 9460 5700 9470 5810
rect 9560 5700 9570 5810
rect 9460 5690 9570 5700
rect 9910 5690 10740 5870
rect 11550 5810 11680 6410
rect 12070 5980 12200 6690
rect 12070 5900 12100 5980
rect 12190 5900 12200 5980
rect 12240 5940 12370 7230
rect 12510 7070 12650 7270
rect 12510 6970 12520 7070
rect 12640 6970 12650 7070
rect 12510 6830 12650 6970
rect 12510 6730 12520 6830
rect 12640 6730 12650 6830
rect 12510 6710 12650 6730
rect 12720 7120 13050 7770
rect 12720 6630 13260 7120
rect 12420 6530 13260 6630
rect 12720 6200 13260 6530
rect 12420 6100 13260 6200
rect 12070 5850 12200 5900
rect 13400 5870 13820 7020
rect 13870 6140 13950 7100
rect 14088 6100 16370 6110
rect 14088 6020 14100 6100
rect 14170 6020 14200 6100
rect 14270 6020 14300 6100
rect 14370 6020 16370 6100
rect 14088 6014 16370 6020
rect 12070 5830 12100 5850
rect 11200 5800 11680 5810
rect 11200 5690 11210 5800
rect 11270 5690 11320 5800
rect 11380 5690 11430 5800
rect 11490 5730 12060 5800
rect 11490 5690 11660 5730
rect 7650 5660 7710 5673
rect 7458 5560 9740 5570
rect 7458 5480 9330 5560
rect 9400 5480 9430 5560
rect 9500 5480 9530 5560
rect 9600 5480 9740 5560
rect 7458 5470 9740 5480
rect 7350 5400 10360 5410
rect 7350 5320 8280 5400
rect 8350 5320 8380 5400
rect 8450 5320 8480 5400
rect 8550 5320 10360 5400
rect 7350 5310 10360 5320
rect 10030 5266 10130 5280
rect 10030 5232 10037 5266
rect 10071 5232 10130 5266
rect 10030 5220 10130 5232
rect 10030 5192 10040 5220
rect 10030 5158 10037 5192
rect 10030 5140 10040 5158
rect 10120 5140 10130 5220
rect 7350 5110 7520 5120
rect 7350 5000 7360 5110
rect 7420 5075 7450 5110
rect 7420 5000 7450 5033
rect 7510 5000 7520 5110
rect 7350 4990 7520 5000
rect 10030 5100 10130 5140
rect 10030 5020 10040 5100
rect 10120 5020 10130 5100
rect 10030 4953 10130 5020
rect 10460 5180 10740 5690
rect 11050 5550 11160 5690
rect 11050 5470 11060 5550
rect 11150 5470 11160 5550
rect 11050 5450 11160 5470
rect 11050 5370 11060 5450
rect 11150 5370 11160 5450
rect 11050 5320 11160 5370
rect 11200 5680 11660 5690
rect 11200 5290 11260 5680
rect 11300 5390 11550 5630
rect 11590 5300 11660 5680
rect 11690 5660 11770 5680
rect 11690 5600 11700 5660
rect 11760 5600 11770 5660
rect 11690 5550 11770 5600
rect 11690 5490 11700 5550
rect 11760 5490 11770 5550
rect 11690 5330 11770 5490
rect 11980 5330 12060 5730
rect 12090 5770 12100 5830
rect 12190 5810 12200 5850
rect 12190 5770 12540 5810
rect 12090 5680 12540 5770
rect 12090 5290 12160 5680
rect 12200 5390 12450 5630
rect 12490 5290 12540 5680
rect 12590 5550 12700 5700
rect 12590 5470 12600 5550
rect 12690 5470 12700 5550
rect 12590 5450 12700 5470
rect 12590 5370 12600 5450
rect 12690 5370 12700 5450
rect 12590 5330 12700 5370
rect 12990 5690 13820 5870
rect 16110 5833 16180 5850
rect 14250 5810 14380 5820
rect 14250 5690 14260 5810
rect 14370 5690 14380 5810
rect 12990 5180 13270 5690
rect 14250 5680 14380 5690
rect 16110 5794 16122 5833
rect 16159 5794 16180 5833
rect 16110 5718 16180 5794
rect 16110 5679 16122 5718
rect 16159 5679 16180 5718
rect 16110 5650 16180 5679
rect 14088 5560 16360 5570
rect 14088 5480 14100 5560
rect 14180 5480 14210 5560
rect 14290 5480 14320 5560
rect 14400 5480 16360 5560
rect 14088 5470 16360 5480
rect 10460 5000 13270 5180
rect 10030 4919 10038 4953
rect 10072 4919 10130 4953
rect 10030 4900 10130 4919
rect 7350 4860 10360 4870
rect 7350 4780 9330 4860
rect 9400 4780 9430 4860
rect 9500 4780 9530 4860
rect 9600 4780 10360 4860
rect 7350 4770 10360 4780
rect 7450 4700 10180 4710
rect 7450 4620 8280 4700
rect 8350 4620 8380 4700
rect 8450 4620 8480 4700
rect 8550 4620 10180 4700
rect 7450 4610 10180 4620
rect 11320 4440 11420 4900
rect 11540 4500 12280 5000
rect 7830 4430 11420 4440
rect 7460 4383 7550 4410
rect 7460 4319 7484 4383
rect 7541 4319 7550 4383
rect 7460 4290 7550 4319
rect 7830 4300 7840 4430
rect 7900 4300 7930 4430
rect 7990 4300 8760 4430
rect 8860 4300 8890 4430
rect 8990 4300 9030 4430
rect 9130 4384 11420 4430
rect 9130 4325 9766 4384
rect 9800 4373 11420 4384
rect 9800 4339 9839 4373
rect 9904 4339 11420 4373
rect 9800 4325 11420 4339
rect 9130 4300 11420 4325
rect 7830 4290 11420 4300
rect 12620 4360 13430 4840
rect 12620 4170 12730 4360
rect 13320 4170 13430 4360
rect 7450 4160 13430 4170
rect 7450 4080 9330 4160
rect 9400 4080 9430 4160
rect 9500 4080 9530 4160
rect 9600 4080 13430 4160
rect 7450 4070 13430 4080
<< via1 >>
rect 10320 8390 10410 8500
rect 10440 8466 10530 8500
rect 10560 8466 10650 8500
rect 10440 8428 10478 8466
rect 10478 8428 10530 8466
rect 10440 8390 10530 8428
rect 10560 8427 10572 8466
rect 10572 8427 10637 8466
rect 10637 8427 10650 8466
rect 10560 8390 10650 8427
rect 10560 8170 10640 8250
rect 10670 8170 10750 8250
rect 10780 8170 10860 8250
rect 8280 6020 8350 6100
rect 8380 6020 8450 6100
rect 8480 6020 8550 6100
rect 9460 6020 9530 6100
rect 9560 6020 9630 6100
rect 9660 6020 9730 6100
rect 11700 7280 11780 7400
rect 11810 7280 11940 7400
rect 11970 7280 12050 7400
rect 11940 7020 12010 7090
rect 11940 6840 12010 6910
rect 11590 6610 11650 6670
rect 11590 6510 11650 6570
rect 11590 6410 11650 6470
rect 9470 5780 9560 5810
rect 9470 5720 9480 5780
rect 9480 5720 9540 5780
rect 9540 5720 9560 5780
rect 9470 5700 9560 5720
rect 12100 5900 12190 5980
rect 14100 6020 14170 6100
rect 14200 6020 14270 6100
rect 14300 6020 14370 6100
rect 11210 5690 11270 5800
rect 11320 5690 11380 5800
rect 11430 5690 11490 5800
rect 9330 5480 9400 5560
rect 9430 5480 9500 5560
rect 9530 5480 9600 5560
rect 8280 5320 8350 5400
rect 8380 5320 8450 5400
rect 8480 5320 8550 5400
rect 10040 5192 10120 5220
rect 10040 5158 10071 5192
rect 10071 5158 10120 5192
rect 10040 5140 10120 5158
rect 7360 5075 7420 5110
rect 7450 5075 7510 5110
rect 7360 5033 7382 5075
rect 7382 5033 7420 5075
rect 7450 5033 7463 5075
rect 7463 5033 7510 5075
rect 7360 5000 7420 5033
rect 7450 5000 7510 5033
rect 10040 5020 10120 5100
rect 11060 5470 11150 5550
rect 11060 5370 11150 5450
rect 11700 5600 11760 5660
rect 11700 5490 11760 5550
rect 12100 5770 12190 5850
rect 12600 5470 12690 5550
rect 12600 5370 12690 5450
rect 14260 5780 14370 5810
rect 14260 5719 14285 5780
rect 14285 5719 14340 5780
rect 14340 5719 14370 5780
rect 14260 5690 14370 5719
rect 14100 5480 14180 5560
rect 14210 5480 14290 5560
rect 14320 5480 14400 5560
rect 9330 4780 9400 4860
rect 9430 4780 9500 4860
rect 9530 4780 9600 4860
rect 8280 4620 8350 4700
rect 8380 4620 8450 4700
rect 8480 4620 8550 4700
rect 7840 4300 7900 4430
rect 7930 4300 7990 4430
rect 8760 4300 8860 4430
rect 8890 4300 8990 4430
rect 9030 4300 9130 4430
rect 9330 4080 9400 4160
rect 9430 4080 9500 4160
rect 9530 4080 9600 4160
<< metal2 >>
rect 8860 8500 10660 8510
rect 8860 8390 10320 8500
rect 10410 8390 10440 8500
rect 10530 8390 10560 8500
rect 10650 8390 10660 8500
rect 8860 8380 10660 8390
rect 8270 6100 8560 6120
rect 8270 6020 8280 6100
rect 8350 6020 8380 6100
rect 8450 6020 8480 6100
rect 8550 6020 8560 6100
rect 8270 5400 8560 6020
rect 8270 5320 8280 5400
rect 8350 5320 8380 5400
rect 8450 5320 8480 5400
rect 8550 5320 8560 5400
rect 7350 5110 8000 5120
rect 7350 5000 7360 5110
rect 7420 5000 7450 5110
rect 7510 5000 8000 5110
rect 7350 4990 8000 5000
rect 7830 4430 8000 4990
rect 8270 4700 8560 5320
rect 8270 4620 8280 4700
rect 8350 4620 8380 4700
rect 8450 4620 8480 4700
rect 8550 4620 8560 4700
rect 8270 4600 8560 4620
rect 8860 4440 9040 8380
rect 9170 8250 10870 8280
rect 9170 8170 10560 8250
rect 10640 8170 10670 8250
rect 10750 8170 10780 8250
rect 10860 8170 10870 8250
rect 9170 8160 10870 8170
rect 9170 5580 9350 8160
rect 11690 7400 12060 7410
rect 11690 7280 11700 7400
rect 11780 7280 11810 7400
rect 11940 7280 11970 7400
rect 12050 7280 12060 7400
rect 11690 7270 12060 7280
rect 11930 7090 12020 7120
rect 11930 7020 11940 7090
rect 12010 7020 12020 7090
rect 11930 6910 12020 7020
rect 11930 6840 11940 6910
rect 12010 6840 12020 6910
rect 11930 6770 12020 6840
rect 11580 6690 12020 6770
rect 11580 6670 11660 6690
rect 11580 6610 11590 6670
rect 11650 6610 11660 6670
rect 11580 6570 11660 6610
rect 11580 6510 11590 6570
rect 11650 6510 11660 6570
rect 11580 6470 11660 6510
rect 11580 6410 11590 6470
rect 11650 6410 11660 6470
rect 11580 6400 11660 6410
rect 9450 6100 9740 6110
rect 9450 6020 9460 6100
rect 9530 6020 9560 6100
rect 9630 6020 9660 6100
rect 9730 6020 9740 6100
rect 9450 6000 9740 6020
rect 14080 6100 14400 6110
rect 14080 6020 14100 6100
rect 14170 6020 14200 6100
rect 14270 6020 14300 6100
rect 14370 6020 14400 6100
rect 14080 6000 14400 6020
rect 12090 5980 12200 5990
rect 12090 5900 12100 5980
rect 12190 5900 12200 5980
rect 12090 5850 12200 5900
rect 9460 5810 11550 5820
rect 12090 5810 12100 5850
rect 9460 5700 9470 5810
rect 9560 5800 11550 5810
rect 9560 5700 11210 5800
rect 9460 5690 11210 5700
rect 11270 5690 11320 5800
rect 11380 5690 11430 5800
rect 11490 5690 11550 5800
rect 9460 5680 11550 5690
rect 11690 5770 12100 5810
rect 12190 5820 12200 5850
rect 12190 5810 14380 5820
rect 12190 5770 14260 5810
rect 11690 5740 14260 5770
rect 11690 5660 11770 5740
rect 12090 5690 14260 5740
rect 14370 5690 14380 5810
rect 12090 5680 14380 5690
rect 11690 5600 11700 5660
rect 11760 5600 11770 5660
rect 9170 5560 9610 5580
rect 9170 5480 9330 5560
rect 9400 5480 9430 5560
rect 9500 5480 9530 5560
rect 9600 5480 9610 5560
rect 9170 5470 9610 5480
rect 9320 4860 9610 5470
rect 11050 5550 11160 5560
rect 11050 5470 11060 5550
rect 11150 5470 11160 5550
rect 11690 5550 11770 5600
rect 14080 5560 14430 5580
rect 11690 5490 11700 5550
rect 11760 5490 11770 5550
rect 11690 5480 11770 5490
rect 12590 5550 12700 5560
rect 11050 5460 11160 5470
rect 10030 5450 11160 5460
rect 12590 5470 12600 5550
rect 12690 5470 12700 5550
rect 14080 5480 14100 5560
rect 14180 5480 14210 5560
rect 14290 5480 14320 5560
rect 14400 5480 14430 5560
rect 14080 5470 14430 5480
rect 12590 5450 12700 5470
rect 10030 5370 11060 5450
rect 11150 5370 12600 5450
rect 12690 5370 12700 5450
rect 10030 5360 12700 5370
rect 10030 5220 10130 5360
rect 10030 5140 10040 5220
rect 10120 5140 10130 5220
rect 10030 5100 10130 5140
rect 10030 5020 10040 5100
rect 10120 5020 10130 5100
rect 10030 5010 10130 5020
rect 9320 4780 9330 4860
rect 9400 4780 9430 4860
rect 9500 4780 9530 4860
rect 9600 4780 9610 4860
rect 7830 4300 7840 4430
rect 7900 4300 7930 4430
rect 7990 4300 8000 4430
rect 7830 4290 8000 4300
rect 8750 4430 9140 4440
rect 8750 4300 8760 4430
rect 8860 4300 8890 4430
rect 8990 4300 9030 4430
rect 9130 4300 9140 4430
rect 8750 4290 9140 4300
rect 9320 4160 9610 4780
rect 9320 4080 9330 4160
rect 9400 4080 9430 4160
rect 9500 4080 9530 4160
rect 9600 4080 9610 4160
rect 9320 4070 9610 4080
<< via2 >>
rect 11700 7280 11780 7400
rect 11810 7280 11940 7400
rect 11970 7280 12050 7400
rect 9460 6020 9530 6100
rect 9560 6020 9630 6100
rect 9660 6020 9730 6100
rect 14100 6020 14170 6100
rect 14200 6020 14270 6100
rect 14300 6020 14370 6100
rect 9330 5480 9400 5560
rect 9430 5480 9500 5560
rect 9530 5480 9600 5560
rect 14100 5480 14180 5560
rect 14210 5480 14290 5560
rect 14320 5480 14400 5560
<< metal3 >>
rect 11690 7400 12060 7410
rect 11690 7280 11700 7400
rect 11780 7280 11810 7400
rect 11940 7280 11970 7400
rect 12050 7280 12060 7400
rect 11690 7270 12060 7280
rect 11810 6110 11940 7270
rect 9450 6100 14400 6110
rect 9450 6020 9460 6100
rect 9530 6020 9560 6100
rect 9630 6020 9660 6100
rect 9730 6020 14100 6100
rect 14170 6020 14200 6100
rect 14270 6020 14300 6100
rect 14370 6020 14400 6100
rect 9450 6000 14400 6020
rect 9320 5560 14430 5580
rect 9170 5480 9330 5560
rect 9400 5480 9430 5560
rect 9500 5480 9530 5560
rect 9600 5480 14100 5560
rect 14180 5480 14210 5560
rect 14290 5480 14320 5560
rect 14400 5480 14430 5560
rect 9170 5470 14430 5480
use sky130_fd_pr__pfet_01v8_FBQ47L  XM1
timestamp 1666924120
transform 0 1 12500 1 0 7901
box -161 -600 169 560
use sky130_fd_pr__pfet_01v8_5AQ4BN  XM2
timestamp 1666923623
transform 0 -1 11220 1 0 7901
box -161 -620 179 560
use sky130_fd_pr__nfet_01v8_ZRN2GS  XM4
timestamp 1667435063
transform 0 -1 10398 -1 0 6609
box -509 -532 509 598
use sky130_fd_pr__nfet_01v8_ZCCU26  XM9
timestamp 1667500205
transform 0 1 12448 -1 0 4669
box -269 -1088 269 1028
use sky130_fd_pr__nfet_01v8_ZZU2YL  XM13
timestamp 1667436771
transform 0 1 11279 -1 0 5511
box -221 -179 221 119
use sky130_fd_pr__nfet_01v8_ZRN2GS  sky130_fd_pr__nfet_01v8_ZRN2GS_0
timestamp 1667435063
transform 0 1 13332 1 0 6609
box -509 -532 509 598
use sky130_fd_pr__nfet_01v8_ZZU2YL  sky130_fd_pr__nfet_01v8_ZZU2YL_0
timestamp 1667436771
transform 0 1 12179 1 0 5511
box -221 -179 221 119
use sky130_fd_pr__nfet_01v8_ZZU2YL  sky130_fd_pr__nfet_01v8_ZZU2YL_1
timestamp 1667436771
transform 0 -1 11569 1 0 5511
box -221 -179 221 119
use sky130_fd_pr__nfet_01v8_ZZU2YL  sky130_fd_pr__nfet_01v8_ZZU2YL_2
timestamp 1667436771
transform 0 -1 12469 1 0 5511
box -221 -179 221 119
use sky130_fd_pr__pfet_01v8_QPTUVJ  sky130_fd_pr__pfet_01v8_QPTUVJ_0
timestamp 1667435677
transform 0 -1 11529 1 0 7007
box -257 -271 263 219
use sky130_fd_pr__pfet_01v8_QPTUVJ  sky130_fd_pr__pfet_01v8_QPTUVJ_1
timestamp 1667435677
transform 0 1 12221 1 0 7007
box -257 -271 263 219
use sky130_fd_pr__pfet_01v8_RPBXXN  sky130_fd_pr__pfet_01v8_RPBXXN_0
timestamp 1666924247
transform 0 -1 12221 -1 0 6249
box -451 -269 449 221
use sky130_fd_pr__pfet_01v8_RPBXXN  sky130_fd_pr__pfet_01v8_RPBXXN_1
timestamp 1666924247
transform 0 1 11529 -1 0 6249
box -451 -269 449 221
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 10268 0 1 4818
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1662439860
transform 1 0 14088 0 1 5518
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1662439860
transform 1 0 9648 0 1 5518
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1662439860
transform 1 0 10088 0 1 4118
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1662439860
transform 1 0 11558 0 1 8208
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  x1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14258 0 1 5518
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14618 0 1 5518
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 15258 0 1 5518
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x4
timestamp 1662439860
transform -1 0 9564 0 1 5518
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x5
timestamp 1662439860
transform -1 0 9200 0 1 5518
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x6
timestamp 1662439860
transform -1 0 8562 0 1 5518
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x7
timestamp 1662439860
transform 1 0 7458 0 1 4118
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 7358 0 1 4818
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9818 0 1 4818
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x10
timestamp 1662439860
transform 1 0 8178 0 1 4818
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8998 0 1 4818
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x12
timestamp 1662439860
transform 1 0 7818 0 1 4118
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  x13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 10558 0 1 8208
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x14
timestamp 1662439860
transform 1 0 8268 0 1 4118
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x15
timestamp 1662439860
transform 1 0 8898 0 1 4118
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  x16
timestamp 1662439860
transform 1 0 10918 0 1 8208
box -38 -48 590 592
<< labels >>
flabel nwell s 8518 6045 8552 6079 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
rlabel metal3 9730 6000 14100 6110 1 VDD
port 5 n
rlabel metal1 9600 4070 13430 4170 1 VSS
port 6 n
rlabel metal1 9780 6120 9860 7080 1 Vin_p
port 7 n
rlabel metal1 7650 5712 7710 5791 1 Out_n
port 8 n
rlabel metal1 13870 6140 13950 7100 1 Vin_n
port 9 n
rlabel metal1 16110 5718 16180 5794 1 Out_p
port 10 n
rlabel metal1 7460 4290 7484 4410 1 ext_clk
port 11 n
<< end >>
