magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< error_p >>
rect -2227 31620 -2167 36030
rect -2147 31620 -2087 36030
rect -1508 31620 -1448 36030
rect -1428 31620 -1368 36030
rect -789 31620 -729 36030
rect -709 31620 -649 36030
rect -70 31620 -10 36030
rect 10 31620 70 36030
rect 649 31620 709 36030
rect 729 31620 789 36030
rect 1368 31620 1428 36030
rect 1448 31620 1508 36030
rect 2087 31620 2147 36030
rect 2167 31620 2227 36030
rect -2227 27110 -2167 31520
rect -2147 27110 -2087 31520
rect -1508 27110 -1448 31520
rect -1428 27110 -1368 31520
rect -789 27110 -729 31520
rect -709 27110 -649 31520
rect -70 27110 -10 31520
rect 10 27110 70 31520
rect 649 27110 709 31520
rect 729 27110 789 31520
rect 1368 27110 1428 31520
rect 1448 27110 1508 31520
rect 2087 27110 2147 31520
rect 2167 27110 2227 31520
rect -2227 22600 -2167 27010
rect -2147 22600 -2087 27010
rect -1508 22600 -1448 27010
rect -1428 22600 -1368 27010
rect -789 22600 -729 27010
rect -709 22600 -649 27010
rect -70 22600 -10 27010
rect 10 22600 70 27010
rect 649 22600 709 27010
rect 729 22600 789 27010
rect 1368 22600 1428 27010
rect 1448 22600 1508 27010
rect 2087 22600 2147 27010
rect 2167 22600 2227 27010
rect -2227 18090 -2167 22500
rect -2147 18090 -2087 22500
rect -1508 18090 -1448 22500
rect -1428 18090 -1368 22500
rect -789 18090 -729 22500
rect -709 18090 -649 22500
rect -70 18090 -10 22500
rect 10 18090 70 22500
rect 649 18090 709 22500
rect 729 18090 789 22500
rect 1368 18090 1428 22500
rect 1448 18090 1508 22500
rect 2087 18090 2147 22500
rect 2167 18090 2227 22500
rect -2227 13580 -2167 17990
rect -2147 13580 -2087 17990
rect -1508 13580 -1448 17990
rect -1428 13580 -1368 17990
rect -789 13580 -729 17990
rect -709 13580 -649 17990
rect -70 13580 -10 17990
rect 10 13580 70 17990
rect 649 13580 709 17990
rect 729 13580 789 17990
rect 1368 13580 1428 17990
rect 1448 13580 1508 17990
rect 2087 13580 2147 17990
rect 2167 13580 2227 17990
rect -2227 9070 -2167 13480
rect -2147 9070 -2087 13480
rect -1508 9070 -1448 13480
rect -1428 9070 -1368 13480
rect -789 9070 -729 13480
rect -709 9070 -649 13480
rect -70 9070 -10 13480
rect 10 9070 70 13480
rect 649 9070 709 13480
rect 729 9070 789 13480
rect 1368 9070 1428 13480
rect 1448 9070 1508 13480
rect 2087 9070 2147 13480
rect 2167 9070 2227 13480
rect -2227 4560 -2167 8970
rect -2147 4560 -2087 8970
rect -1508 4560 -1448 8970
rect -1428 4560 -1368 8970
rect -789 4560 -729 8970
rect -709 4560 -649 8970
rect -70 4560 -10 8970
rect 10 4560 70 8970
rect 649 4560 709 8970
rect 729 4560 789 8970
rect 1368 4560 1428 8970
rect 1448 4560 1508 8970
rect 2087 4560 2147 8970
rect 2167 4560 2227 8970
rect -2227 50 -2167 4460
rect -2147 50 -2087 4460
rect -1508 50 -1448 4460
rect -1428 50 -1368 4460
rect -789 50 -729 4460
rect -709 50 -649 4460
rect -70 50 -10 4460
rect 10 50 70 4460
rect 649 50 709 4460
rect 729 50 789 4460
rect 1368 50 1428 4460
rect 1448 50 1508 4460
rect 2087 50 2147 4460
rect 2167 50 2227 4460
rect -2227 -4460 -2167 -50
rect -2147 -4460 -2087 -50
rect -1508 -4460 -1448 -50
rect -1428 -4460 -1368 -50
rect -789 -4460 -729 -50
rect -709 -4460 -649 -50
rect -70 -4460 -10 -50
rect 10 -4460 70 -50
rect 649 -4460 709 -50
rect 729 -4460 789 -50
rect 1368 -4460 1428 -50
rect 1448 -4460 1508 -50
rect 2087 -4460 2147 -50
rect 2167 -4460 2227 -50
rect -2227 -8970 -2167 -4560
rect -2147 -8970 -2087 -4560
rect -1508 -8970 -1448 -4560
rect -1428 -8970 -1368 -4560
rect -789 -8970 -729 -4560
rect -709 -8970 -649 -4560
rect -70 -8970 -10 -4560
rect 10 -8970 70 -4560
rect 649 -8970 709 -4560
rect 729 -8970 789 -4560
rect 1368 -8970 1428 -4560
rect 1448 -8970 1508 -4560
rect 2087 -8970 2147 -4560
rect 2167 -8970 2227 -4560
rect -2227 -13480 -2167 -9070
rect -2147 -13480 -2087 -9070
rect -1508 -13480 -1448 -9070
rect -1428 -13480 -1368 -9070
rect -789 -13480 -729 -9070
rect -709 -13480 -649 -9070
rect -70 -13480 -10 -9070
rect 10 -13480 70 -9070
rect 649 -13480 709 -9070
rect 729 -13480 789 -9070
rect 1368 -13480 1428 -9070
rect 1448 -13480 1508 -9070
rect 2087 -13480 2147 -9070
rect 2167 -13480 2227 -9070
rect -2227 -17990 -2167 -13580
rect -2147 -17990 -2087 -13580
rect -1508 -17990 -1448 -13580
rect -1428 -17990 -1368 -13580
rect -789 -17990 -729 -13580
rect -709 -17990 -649 -13580
rect -70 -17990 -10 -13580
rect 10 -17990 70 -13580
rect 649 -17990 709 -13580
rect 729 -17990 789 -13580
rect 1368 -17990 1428 -13580
rect 1448 -17990 1508 -13580
rect 2087 -17990 2147 -13580
rect 2167 -17990 2227 -13580
rect -2227 -22500 -2167 -18090
rect -2147 -22500 -2087 -18090
rect -1508 -22500 -1448 -18090
rect -1428 -22500 -1368 -18090
rect -789 -22500 -729 -18090
rect -709 -22500 -649 -18090
rect -70 -22500 -10 -18090
rect 10 -22500 70 -18090
rect 649 -22500 709 -18090
rect 729 -22500 789 -18090
rect 1368 -22500 1428 -18090
rect 1448 -22500 1508 -18090
rect 2087 -22500 2147 -18090
rect 2167 -22500 2227 -18090
rect -2227 -27010 -2167 -22600
rect -2147 -27010 -2087 -22600
rect -1508 -27010 -1448 -22600
rect -1428 -27010 -1368 -22600
rect -789 -27010 -729 -22600
rect -709 -27010 -649 -22600
rect -70 -27010 -10 -22600
rect 10 -27010 70 -22600
rect 649 -27010 709 -22600
rect 729 -27010 789 -22600
rect 1368 -27010 1428 -22600
rect 1448 -27010 1508 -22600
rect 2087 -27010 2147 -22600
rect 2167 -27010 2227 -22600
rect -2227 -31520 -2167 -27110
rect -2147 -31520 -2087 -27110
rect -1508 -31520 -1448 -27110
rect -1428 -31520 -1368 -27110
rect -789 -31520 -729 -27110
rect -709 -31520 -649 -27110
rect -70 -31520 -10 -27110
rect 10 -31520 70 -27110
rect 649 -31520 709 -27110
rect 729 -31520 789 -27110
rect 1368 -31520 1428 -27110
rect 1448 -31520 1508 -27110
rect 2087 -31520 2147 -27110
rect 2167 -31520 2227 -27110
rect -2227 -36030 -2167 -31620
rect -2147 -36030 -2087 -31620
rect -1508 -36030 -1448 -31620
rect -1428 -36030 -1368 -31620
rect -789 -36030 -729 -31620
rect -709 -36030 -649 -31620
rect -70 -36030 -10 -31620
rect 10 -36030 70 -31620
rect 649 -36030 709 -31620
rect 729 -36030 789 -31620
rect 1368 -36030 1428 -31620
rect 1448 -36030 1508 -31620
rect 2087 -36030 2147 -31620
rect 2167 -36030 2227 -31620
<< metal3 >>
rect -2866 36002 -2167 36030
rect -2866 31648 -2251 36002
rect -2187 31648 -2167 36002
rect -2866 31620 -2167 31648
rect -2147 36002 -1448 36030
rect -2147 31648 -1532 36002
rect -1468 31648 -1448 36002
rect -2147 31620 -1448 31648
rect -1428 36002 -729 36030
rect -1428 31648 -813 36002
rect -749 31648 -729 36002
rect -1428 31620 -729 31648
rect -709 36002 -10 36030
rect -709 31648 -94 36002
rect -30 31648 -10 36002
rect -709 31620 -10 31648
rect 10 36002 709 36030
rect 10 31648 625 36002
rect 689 31648 709 36002
rect 10 31620 709 31648
rect 729 36002 1428 36030
rect 729 31648 1344 36002
rect 1408 31648 1428 36002
rect 729 31620 1428 31648
rect 1448 36002 2147 36030
rect 1448 31648 2063 36002
rect 2127 31648 2147 36002
rect 1448 31620 2147 31648
rect 2167 36002 2866 36030
rect 2167 31648 2782 36002
rect 2846 31648 2866 36002
rect 2167 31620 2866 31648
rect -2866 31492 -2167 31520
rect -2866 27138 -2251 31492
rect -2187 27138 -2167 31492
rect -2866 27110 -2167 27138
rect -2147 31492 -1448 31520
rect -2147 27138 -1532 31492
rect -1468 27138 -1448 31492
rect -2147 27110 -1448 27138
rect -1428 31492 -729 31520
rect -1428 27138 -813 31492
rect -749 27138 -729 31492
rect -1428 27110 -729 27138
rect -709 31492 -10 31520
rect -709 27138 -94 31492
rect -30 27138 -10 31492
rect -709 27110 -10 27138
rect 10 31492 709 31520
rect 10 27138 625 31492
rect 689 27138 709 31492
rect 10 27110 709 27138
rect 729 31492 1428 31520
rect 729 27138 1344 31492
rect 1408 27138 1428 31492
rect 729 27110 1428 27138
rect 1448 31492 2147 31520
rect 1448 27138 2063 31492
rect 2127 27138 2147 31492
rect 1448 27110 2147 27138
rect 2167 31492 2866 31520
rect 2167 27138 2782 31492
rect 2846 27138 2866 31492
rect 2167 27110 2866 27138
rect -2866 26982 -2167 27010
rect -2866 22628 -2251 26982
rect -2187 22628 -2167 26982
rect -2866 22600 -2167 22628
rect -2147 26982 -1448 27010
rect -2147 22628 -1532 26982
rect -1468 22628 -1448 26982
rect -2147 22600 -1448 22628
rect -1428 26982 -729 27010
rect -1428 22628 -813 26982
rect -749 22628 -729 26982
rect -1428 22600 -729 22628
rect -709 26982 -10 27010
rect -709 22628 -94 26982
rect -30 22628 -10 26982
rect -709 22600 -10 22628
rect 10 26982 709 27010
rect 10 22628 625 26982
rect 689 22628 709 26982
rect 10 22600 709 22628
rect 729 26982 1428 27010
rect 729 22628 1344 26982
rect 1408 22628 1428 26982
rect 729 22600 1428 22628
rect 1448 26982 2147 27010
rect 1448 22628 2063 26982
rect 2127 22628 2147 26982
rect 1448 22600 2147 22628
rect 2167 26982 2866 27010
rect 2167 22628 2782 26982
rect 2846 22628 2866 26982
rect 2167 22600 2866 22628
rect -2866 22472 -2167 22500
rect -2866 18118 -2251 22472
rect -2187 18118 -2167 22472
rect -2866 18090 -2167 18118
rect -2147 22472 -1448 22500
rect -2147 18118 -1532 22472
rect -1468 18118 -1448 22472
rect -2147 18090 -1448 18118
rect -1428 22472 -729 22500
rect -1428 18118 -813 22472
rect -749 18118 -729 22472
rect -1428 18090 -729 18118
rect -709 22472 -10 22500
rect -709 18118 -94 22472
rect -30 18118 -10 22472
rect -709 18090 -10 18118
rect 10 22472 709 22500
rect 10 18118 625 22472
rect 689 18118 709 22472
rect 10 18090 709 18118
rect 729 22472 1428 22500
rect 729 18118 1344 22472
rect 1408 18118 1428 22472
rect 729 18090 1428 18118
rect 1448 22472 2147 22500
rect 1448 18118 2063 22472
rect 2127 18118 2147 22472
rect 1448 18090 2147 18118
rect 2167 22472 2866 22500
rect 2167 18118 2782 22472
rect 2846 18118 2866 22472
rect 2167 18090 2866 18118
rect -2866 17962 -2167 17990
rect -2866 13608 -2251 17962
rect -2187 13608 -2167 17962
rect -2866 13580 -2167 13608
rect -2147 17962 -1448 17990
rect -2147 13608 -1532 17962
rect -1468 13608 -1448 17962
rect -2147 13580 -1448 13608
rect -1428 17962 -729 17990
rect -1428 13608 -813 17962
rect -749 13608 -729 17962
rect -1428 13580 -729 13608
rect -709 17962 -10 17990
rect -709 13608 -94 17962
rect -30 13608 -10 17962
rect -709 13580 -10 13608
rect 10 17962 709 17990
rect 10 13608 625 17962
rect 689 13608 709 17962
rect 10 13580 709 13608
rect 729 17962 1428 17990
rect 729 13608 1344 17962
rect 1408 13608 1428 17962
rect 729 13580 1428 13608
rect 1448 17962 2147 17990
rect 1448 13608 2063 17962
rect 2127 13608 2147 17962
rect 1448 13580 2147 13608
rect 2167 17962 2866 17990
rect 2167 13608 2782 17962
rect 2846 13608 2866 17962
rect 2167 13580 2866 13608
rect -2866 13452 -2167 13480
rect -2866 9098 -2251 13452
rect -2187 9098 -2167 13452
rect -2866 9070 -2167 9098
rect -2147 13452 -1448 13480
rect -2147 9098 -1532 13452
rect -1468 9098 -1448 13452
rect -2147 9070 -1448 9098
rect -1428 13452 -729 13480
rect -1428 9098 -813 13452
rect -749 9098 -729 13452
rect -1428 9070 -729 9098
rect -709 13452 -10 13480
rect -709 9098 -94 13452
rect -30 9098 -10 13452
rect -709 9070 -10 9098
rect 10 13452 709 13480
rect 10 9098 625 13452
rect 689 9098 709 13452
rect 10 9070 709 9098
rect 729 13452 1428 13480
rect 729 9098 1344 13452
rect 1408 9098 1428 13452
rect 729 9070 1428 9098
rect 1448 13452 2147 13480
rect 1448 9098 2063 13452
rect 2127 9098 2147 13452
rect 1448 9070 2147 9098
rect 2167 13452 2866 13480
rect 2167 9098 2782 13452
rect 2846 9098 2866 13452
rect 2167 9070 2866 9098
rect -2866 8942 -2167 8970
rect -2866 4588 -2251 8942
rect -2187 4588 -2167 8942
rect -2866 4560 -2167 4588
rect -2147 8942 -1448 8970
rect -2147 4588 -1532 8942
rect -1468 4588 -1448 8942
rect -2147 4560 -1448 4588
rect -1428 8942 -729 8970
rect -1428 4588 -813 8942
rect -749 4588 -729 8942
rect -1428 4560 -729 4588
rect -709 8942 -10 8970
rect -709 4588 -94 8942
rect -30 4588 -10 8942
rect -709 4560 -10 4588
rect 10 8942 709 8970
rect 10 4588 625 8942
rect 689 4588 709 8942
rect 10 4560 709 4588
rect 729 8942 1428 8970
rect 729 4588 1344 8942
rect 1408 4588 1428 8942
rect 729 4560 1428 4588
rect 1448 8942 2147 8970
rect 1448 4588 2063 8942
rect 2127 4588 2147 8942
rect 1448 4560 2147 4588
rect 2167 8942 2866 8970
rect 2167 4588 2782 8942
rect 2846 4588 2866 8942
rect 2167 4560 2866 4588
rect -2866 4432 -2167 4460
rect -2866 78 -2251 4432
rect -2187 78 -2167 4432
rect -2866 50 -2167 78
rect -2147 4432 -1448 4460
rect -2147 78 -1532 4432
rect -1468 78 -1448 4432
rect -2147 50 -1448 78
rect -1428 4432 -729 4460
rect -1428 78 -813 4432
rect -749 78 -729 4432
rect -1428 50 -729 78
rect -709 4432 -10 4460
rect -709 78 -94 4432
rect -30 78 -10 4432
rect -709 50 -10 78
rect 10 4432 709 4460
rect 10 78 625 4432
rect 689 78 709 4432
rect 10 50 709 78
rect 729 4432 1428 4460
rect 729 78 1344 4432
rect 1408 78 1428 4432
rect 729 50 1428 78
rect 1448 4432 2147 4460
rect 1448 78 2063 4432
rect 2127 78 2147 4432
rect 1448 50 2147 78
rect 2167 4432 2866 4460
rect 2167 78 2782 4432
rect 2846 78 2866 4432
rect 2167 50 2866 78
rect -2866 -78 -2167 -50
rect -2866 -4432 -2251 -78
rect -2187 -4432 -2167 -78
rect -2866 -4460 -2167 -4432
rect -2147 -78 -1448 -50
rect -2147 -4432 -1532 -78
rect -1468 -4432 -1448 -78
rect -2147 -4460 -1448 -4432
rect -1428 -78 -729 -50
rect -1428 -4432 -813 -78
rect -749 -4432 -729 -78
rect -1428 -4460 -729 -4432
rect -709 -78 -10 -50
rect -709 -4432 -94 -78
rect -30 -4432 -10 -78
rect -709 -4460 -10 -4432
rect 10 -78 709 -50
rect 10 -4432 625 -78
rect 689 -4432 709 -78
rect 10 -4460 709 -4432
rect 729 -78 1428 -50
rect 729 -4432 1344 -78
rect 1408 -4432 1428 -78
rect 729 -4460 1428 -4432
rect 1448 -78 2147 -50
rect 1448 -4432 2063 -78
rect 2127 -4432 2147 -78
rect 1448 -4460 2147 -4432
rect 2167 -78 2866 -50
rect 2167 -4432 2782 -78
rect 2846 -4432 2866 -78
rect 2167 -4460 2866 -4432
rect -2866 -4588 -2167 -4560
rect -2866 -8942 -2251 -4588
rect -2187 -8942 -2167 -4588
rect -2866 -8970 -2167 -8942
rect -2147 -4588 -1448 -4560
rect -2147 -8942 -1532 -4588
rect -1468 -8942 -1448 -4588
rect -2147 -8970 -1448 -8942
rect -1428 -4588 -729 -4560
rect -1428 -8942 -813 -4588
rect -749 -8942 -729 -4588
rect -1428 -8970 -729 -8942
rect -709 -4588 -10 -4560
rect -709 -8942 -94 -4588
rect -30 -8942 -10 -4588
rect -709 -8970 -10 -8942
rect 10 -4588 709 -4560
rect 10 -8942 625 -4588
rect 689 -8942 709 -4588
rect 10 -8970 709 -8942
rect 729 -4588 1428 -4560
rect 729 -8942 1344 -4588
rect 1408 -8942 1428 -4588
rect 729 -8970 1428 -8942
rect 1448 -4588 2147 -4560
rect 1448 -8942 2063 -4588
rect 2127 -8942 2147 -4588
rect 1448 -8970 2147 -8942
rect 2167 -4588 2866 -4560
rect 2167 -8942 2782 -4588
rect 2846 -8942 2866 -4588
rect 2167 -8970 2866 -8942
rect -2866 -9098 -2167 -9070
rect -2866 -13452 -2251 -9098
rect -2187 -13452 -2167 -9098
rect -2866 -13480 -2167 -13452
rect -2147 -9098 -1448 -9070
rect -2147 -13452 -1532 -9098
rect -1468 -13452 -1448 -9098
rect -2147 -13480 -1448 -13452
rect -1428 -9098 -729 -9070
rect -1428 -13452 -813 -9098
rect -749 -13452 -729 -9098
rect -1428 -13480 -729 -13452
rect -709 -9098 -10 -9070
rect -709 -13452 -94 -9098
rect -30 -13452 -10 -9098
rect -709 -13480 -10 -13452
rect 10 -9098 709 -9070
rect 10 -13452 625 -9098
rect 689 -13452 709 -9098
rect 10 -13480 709 -13452
rect 729 -9098 1428 -9070
rect 729 -13452 1344 -9098
rect 1408 -13452 1428 -9098
rect 729 -13480 1428 -13452
rect 1448 -9098 2147 -9070
rect 1448 -13452 2063 -9098
rect 2127 -13452 2147 -9098
rect 1448 -13480 2147 -13452
rect 2167 -9098 2866 -9070
rect 2167 -13452 2782 -9098
rect 2846 -13452 2866 -9098
rect 2167 -13480 2866 -13452
rect -2866 -13608 -2167 -13580
rect -2866 -17962 -2251 -13608
rect -2187 -17962 -2167 -13608
rect -2866 -17990 -2167 -17962
rect -2147 -13608 -1448 -13580
rect -2147 -17962 -1532 -13608
rect -1468 -17962 -1448 -13608
rect -2147 -17990 -1448 -17962
rect -1428 -13608 -729 -13580
rect -1428 -17962 -813 -13608
rect -749 -17962 -729 -13608
rect -1428 -17990 -729 -17962
rect -709 -13608 -10 -13580
rect -709 -17962 -94 -13608
rect -30 -17962 -10 -13608
rect -709 -17990 -10 -17962
rect 10 -13608 709 -13580
rect 10 -17962 625 -13608
rect 689 -17962 709 -13608
rect 10 -17990 709 -17962
rect 729 -13608 1428 -13580
rect 729 -17962 1344 -13608
rect 1408 -17962 1428 -13608
rect 729 -17990 1428 -17962
rect 1448 -13608 2147 -13580
rect 1448 -17962 2063 -13608
rect 2127 -17962 2147 -13608
rect 1448 -17990 2147 -17962
rect 2167 -13608 2866 -13580
rect 2167 -17962 2782 -13608
rect 2846 -17962 2866 -13608
rect 2167 -17990 2866 -17962
rect -2866 -18118 -2167 -18090
rect -2866 -22472 -2251 -18118
rect -2187 -22472 -2167 -18118
rect -2866 -22500 -2167 -22472
rect -2147 -18118 -1448 -18090
rect -2147 -22472 -1532 -18118
rect -1468 -22472 -1448 -18118
rect -2147 -22500 -1448 -22472
rect -1428 -18118 -729 -18090
rect -1428 -22472 -813 -18118
rect -749 -22472 -729 -18118
rect -1428 -22500 -729 -22472
rect -709 -18118 -10 -18090
rect -709 -22472 -94 -18118
rect -30 -22472 -10 -18118
rect -709 -22500 -10 -22472
rect 10 -18118 709 -18090
rect 10 -22472 625 -18118
rect 689 -22472 709 -18118
rect 10 -22500 709 -22472
rect 729 -18118 1428 -18090
rect 729 -22472 1344 -18118
rect 1408 -22472 1428 -18118
rect 729 -22500 1428 -22472
rect 1448 -18118 2147 -18090
rect 1448 -22472 2063 -18118
rect 2127 -22472 2147 -18118
rect 1448 -22500 2147 -22472
rect 2167 -18118 2866 -18090
rect 2167 -22472 2782 -18118
rect 2846 -22472 2866 -18118
rect 2167 -22500 2866 -22472
rect -2866 -22628 -2167 -22600
rect -2866 -26982 -2251 -22628
rect -2187 -26982 -2167 -22628
rect -2866 -27010 -2167 -26982
rect -2147 -22628 -1448 -22600
rect -2147 -26982 -1532 -22628
rect -1468 -26982 -1448 -22628
rect -2147 -27010 -1448 -26982
rect -1428 -22628 -729 -22600
rect -1428 -26982 -813 -22628
rect -749 -26982 -729 -22628
rect -1428 -27010 -729 -26982
rect -709 -22628 -10 -22600
rect -709 -26982 -94 -22628
rect -30 -26982 -10 -22628
rect -709 -27010 -10 -26982
rect 10 -22628 709 -22600
rect 10 -26982 625 -22628
rect 689 -26982 709 -22628
rect 10 -27010 709 -26982
rect 729 -22628 1428 -22600
rect 729 -26982 1344 -22628
rect 1408 -26982 1428 -22628
rect 729 -27010 1428 -26982
rect 1448 -22628 2147 -22600
rect 1448 -26982 2063 -22628
rect 2127 -26982 2147 -22628
rect 1448 -27010 2147 -26982
rect 2167 -22628 2866 -22600
rect 2167 -26982 2782 -22628
rect 2846 -26982 2866 -22628
rect 2167 -27010 2866 -26982
rect -2866 -27138 -2167 -27110
rect -2866 -31492 -2251 -27138
rect -2187 -31492 -2167 -27138
rect -2866 -31520 -2167 -31492
rect -2147 -27138 -1448 -27110
rect -2147 -31492 -1532 -27138
rect -1468 -31492 -1448 -27138
rect -2147 -31520 -1448 -31492
rect -1428 -27138 -729 -27110
rect -1428 -31492 -813 -27138
rect -749 -31492 -729 -27138
rect -1428 -31520 -729 -31492
rect -709 -27138 -10 -27110
rect -709 -31492 -94 -27138
rect -30 -31492 -10 -27138
rect -709 -31520 -10 -31492
rect 10 -27138 709 -27110
rect 10 -31492 625 -27138
rect 689 -31492 709 -27138
rect 10 -31520 709 -31492
rect 729 -27138 1428 -27110
rect 729 -31492 1344 -27138
rect 1408 -31492 1428 -27138
rect 729 -31520 1428 -31492
rect 1448 -27138 2147 -27110
rect 1448 -31492 2063 -27138
rect 2127 -31492 2147 -27138
rect 1448 -31520 2147 -31492
rect 2167 -27138 2866 -27110
rect 2167 -31492 2782 -27138
rect 2846 -31492 2866 -27138
rect 2167 -31520 2866 -31492
rect -2866 -31648 -2167 -31620
rect -2866 -36002 -2251 -31648
rect -2187 -36002 -2167 -31648
rect -2866 -36030 -2167 -36002
rect -2147 -31648 -1448 -31620
rect -2147 -36002 -1532 -31648
rect -1468 -36002 -1448 -31648
rect -2147 -36030 -1448 -36002
rect -1428 -31648 -729 -31620
rect -1428 -36002 -813 -31648
rect -749 -36002 -729 -31648
rect -1428 -36030 -729 -36002
rect -709 -31648 -10 -31620
rect -709 -36002 -94 -31648
rect -30 -36002 -10 -31648
rect -709 -36030 -10 -36002
rect 10 -31648 709 -31620
rect 10 -36002 625 -31648
rect 689 -36002 709 -31648
rect 10 -36030 709 -36002
rect 729 -31648 1428 -31620
rect 729 -36002 1344 -31648
rect 1408 -36002 1428 -31648
rect 729 -36030 1428 -36002
rect 1448 -31648 2147 -31620
rect 1448 -36002 2063 -31648
rect 2127 -36002 2147 -31648
rect 1448 -36030 2147 -36002
rect 2167 -31648 2866 -31620
rect 2167 -36002 2782 -31648
rect 2846 -36002 2866 -31648
rect 2167 -36030 2866 -36002
<< via3 >>
rect -2251 31648 -2187 36002
rect -1532 31648 -1468 36002
rect -813 31648 -749 36002
rect -94 31648 -30 36002
rect 625 31648 689 36002
rect 1344 31648 1408 36002
rect 2063 31648 2127 36002
rect 2782 31648 2846 36002
rect -2251 27138 -2187 31492
rect -1532 27138 -1468 31492
rect -813 27138 -749 31492
rect -94 27138 -30 31492
rect 625 27138 689 31492
rect 1344 27138 1408 31492
rect 2063 27138 2127 31492
rect 2782 27138 2846 31492
rect -2251 22628 -2187 26982
rect -1532 22628 -1468 26982
rect -813 22628 -749 26982
rect -94 22628 -30 26982
rect 625 22628 689 26982
rect 1344 22628 1408 26982
rect 2063 22628 2127 26982
rect 2782 22628 2846 26982
rect -2251 18118 -2187 22472
rect -1532 18118 -1468 22472
rect -813 18118 -749 22472
rect -94 18118 -30 22472
rect 625 18118 689 22472
rect 1344 18118 1408 22472
rect 2063 18118 2127 22472
rect 2782 18118 2846 22472
rect -2251 13608 -2187 17962
rect -1532 13608 -1468 17962
rect -813 13608 -749 17962
rect -94 13608 -30 17962
rect 625 13608 689 17962
rect 1344 13608 1408 17962
rect 2063 13608 2127 17962
rect 2782 13608 2846 17962
rect -2251 9098 -2187 13452
rect -1532 9098 -1468 13452
rect -813 9098 -749 13452
rect -94 9098 -30 13452
rect 625 9098 689 13452
rect 1344 9098 1408 13452
rect 2063 9098 2127 13452
rect 2782 9098 2846 13452
rect -2251 4588 -2187 8942
rect -1532 4588 -1468 8942
rect -813 4588 -749 8942
rect -94 4588 -30 8942
rect 625 4588 689 8942
rect 1344 4588 1408 8942
rect 2063 4588 2127 8942
rect 2782 4588 2846 8942
rect -2251 78 -2187 4432
rect -1532 78 -1468 4432
rect -813 78 -749 4432
rect -94 78 -30 4432
rect 625 78 689 4432
rect 1344 78 1408 4432
rect 2063 78 2127 4432
rect 2782 78 2846 4432
rect -2251 -4432 -2187 -78
rect -1532 -4432 -1468 -78
rect -813 -4432 -749 -78
rect -94 -4432 -30 -78
rect 625 -4432 689 -78
rect 1344 -4432 1408 -78
rect 2063 -4432 2127 -78
rect 2782 -4432 2846 -78
rect -2251 -8942 -2187 -4588
rect -1532 -8942 -1468 -4588
rect -813 -8942 -749 -4588
rect -94 -8942 -30 -4588
rect 625 -8942 689 -4588
rect 1344 -8942 1408 -4588
rect 2063 -8942 2127 -4588
rect 2782 -8942 2846 -4588
rect -2251 -13452 -2187 -9098
rect -1532 -13452 -1468 -9098
rect -813 -13452 -749 -9098
rect -94 -13452 -30 -9098
rect 625 -13452 689 -9098
rect 1344 -13452 1408 -9098
rect 2063 -13452 2127 -9098
rect 2782 -13452 2846 -9098
rect -2251 -17962 -2187 -13608
rect -1532 -17962 -1468 -13608
rect -813 -17962 -749 -13608
rect -94 -17962 -30 -13608
rect 625 -17962 689 -13608
rect 1344 -17962 1408 -13608
rect 2063 -17962 2127 -13608
rect 2782 -17962 2846 -13608
rect -2251 -22472 -2187 -18118
rect -1532 -22472 -1468 -18118
rect -813 -22472 -749 -18118
rect -94 -22472 -30 -18118
rect 625 -22472 689 -18118
rect 1344 -22472 1408 -18118
rect 2063 -22472 2127 -18118
rect 2782 -22472 2846 -18118
rect -2251 -26982 -2187 -22628
rect -1532 -26982 -1468 -22628
rect -813 -26982 -749 -22628
rect -94 -26982 -30 -22628
rect 625 -26982 689 -22628
rect 1344 -26982 1408 -22628
rect 2063 -26982 2127 -22628
rect 2782 -26982 2846 -22628
rect -2251 -31492 -2187 -27138
rect -1532 -31492 -1468 -27138
rect -813 -31492 -749 -27138
rect -94 -31492 -30 -27138
rect 625 -31492 689 -27138
rect 1344 -31492 1408 -27138
rect 2063 -31492 2127 -27138
rect 2782 -31492 2846 -27138
rect -2251 -36002 -2187 -31648
rect -1532 -36002 -1468 -31648
rect -813 -36002 -749 -31648
rect -94 -36002 -30 -31648
rect 625 -36002 689 -31648
rect 1344 -36002 1408 -31648
rect 2063 -36002 2127 -31648
rect 2782 -36002 2846 -31648
<< mimcap >>
rect -2766 35890 -2366 35930
rect -2766 31760 -2726 35890
rect -2406 31760 -2366 35890
rect -2766 31720 -2366 31760
rect -2047 35890 -1647 35930
rect -2047 31760 -2007 35890
rect -1687 31760 -1647 35890
rect -2047 31720 -1647 31760
rect -1328 35890 -928 35930
rect -1328 31760 -1288 35890
rect -968 31760 -928 35890
rect -1328 31720 -928 31760
rect -609 35890 -209 35930
rect -609 31760 -569 35890
rect -249 31760 -209 35890
rect -609 31720 -209 31760
rect 110 35890 510 35930
rect 110 31760 150 35890
rect 470 31760 510 35890
rect 110 31720 510 31760
rect 829 35890 1229 35930
rect 829 31760 869 35890
rect 1189 31760 1229 35890
rect 829 31720 1229 31760
rect 1548 35890 1948 35930
rect 1548 31760 1588 35890
rect 1908 31760 1948 35890
rect 1548 31720 1948 31760
rect 2267 35890 2667 35930
rect 2267 31760 2307 35890
rect 2627 31760 2667 35890
rect 2267 31720 2667 31760
rect -2766 31380 -2366 31420
rect -2766 27250 -2726 31380
rect -2406 27250 -2366 31380
rect -2766 27210 -2366 27250
rect -2047 31380 -1647 31420
rect -2047 27250 -2007 31380
rect -1687 27250 -1647 31380
rect -2047 27210 -1647 27250
rect -1328 31380 -928 31420
rect -1328 27250 -1288 31380
rect -968 27250 -928 31380
rect -1328 27210 -928 27250
rect -609 31380 -209 31420
rect -609 27250 -569 31380
rect -249 27250 -209 31380
rect -609 27210 -209 27250
rect 110 31380 510 31420
rect 110 27250 150 31380
rect 470 27250 510 31380
rect 110 27210 510 27250
rect 829 31380 1229 31420
rect 829 27250 869 31380
rect 1189 27250 1229 31380
rect 829 27210 1229 27250
rect 1548 31380 1948 31420
rect 1548 27250 1588 31380
rect 1908 27250 1948 31380
rect 1548 27210 1948 27250
rect 2267 31380 2667 31420
rect 2267 27250 2307 31380
rect 2627 27250 2667 31380
rect 2267 27210 2667 27250
rect -2766 26870 -2366 26910
rect -2766 22740 -2726 26870
rect -2406 22740 -2366 26870
rect -2766 22700 -2366 22740
rect -2047 26870 -1647 26910
rect -2047 22740 -2007 26870
rect -1687 22740 -1647 26870
rect -2047 22700 -1647 22740
rect -1328 26870 -928 26910
rect -1328 22740 -1288 26870
rect -968 22740 -928 26870
rect -1328 22700 -928 22740
rect -609 26870 -209 26910
rect -609 22740 -569 26870
rect -249 22740 -209 26870
rect -609 22700 -209 22740
rect 110 26870 510 26910
rect 110 22740 150 26870
rect 470 22740 510 26870
rect 110 22700 510 22740
rect 829 26870 1229 26910
rect 829 22740 869 26870
rect 1189 22740 1229 26870
rect 829 22700 1229 22740
rect 1548 26870 1948 26910
rect 1548 22740 1588 26870
rect 1908 22740 1948 26870
rect 1548 22700 1948 22740
rect 2267 26870 2667 26910
rect 2267 22740 2307 26870
rect 2627 22740 2667 26870
rect 2267 22700 2667 22740
rect -2766 22360 -2366 22400
rect -2766 18230 -2726 22360
rect -2406 18230 -2366 22360
rect -2766 18190 -2366 18230
rect -2047 22360 -1647 22400
rect -2047 18230 -2007 22360
rect -1687 18230 -1647 22360
rect -2047 18190 -1647 18230
rect -1328 22360 -928 22400
rect -1328 18230 -1288 22360
rect -968 18230 -928 22360
rect -1328 18190 -928 18230
rect -609 22360 -209 22400
rect -609 18230 -569 22360
rect -249 18230 -209 22360
rect -609 18190 -209 18230
rect 110 22360 510 22400
rect 110 18230 150 22360
rect 470 18230 510 22360
rect 110 18190 510 18230
rect 829 22360 1229 22400
rect 829 18230 869 22360
rect 1189 18230 1229 22360
rect 829 18190 1229 18230
rect 1548 22360 1948 22400
rect 1548 18230 1588 22360
rect 1908 18230 1948 22360
rect 1548 18190 1948 18230
rect 2267 22360 2667 22400
rect 2267 18230 2307 22360
rect 2627 18230 2667 22360
rect 2267 18190 2667 18230
rect -2766 17850 -2366 17890
rect -2766 13720 -2726 17850
rect -2406 13720 -2366 17850
rect -2766 13680 -2366 13720
rect -2047 17850 -1647 17890
rect -2047 13720 -2007 17850
rect -1687 13720 -1647 17850
rect -2047 13680 -1647 13720
rect -1328 17850 -928 17890
rect -1328 13720 -1288 17850
rect -968 13720 -928 17850
rect -1328 13680 -928 13720
rect -609 17850 -209 17890
rect -609 13720 -569 17850
rect -249 13720 -209 17850
rect -609 13680 -209 13720
rect 110 17850 510 17890
rect 110 13720 150 17850
rect 470 13720 510 17850
rect 110 13680 510 13720
rect 829 17850 1229 17890
rect 829 13720 869 17850
rect 1189 13720 1229 17850
rect 829 13680 1229 13720
rect 1548 17850 1948 17890
rect 1548 13720 1588 17850
rect 1908 13720 1948 17850
rect 1548 13680 1948 13720
rect 2267 17850 2667 17890
rect 2267 13720 2307 17850
rect 2627 13720 2667 17850
rect 2267 13680 2667 13720
rect -2766 13340 -2366 13380
rect -2766 9210 -2726 13340
rect -2406 9210 -2366 13340
rect -2766 9170 -2366 9210
rect -2047 13340 -1647 13380
rect -2047 9210 -2007 13340
rect -1687 9210 -1647 13340
rect -2047 9170 -1647 9210
rect -1328 13340 -928 13380
rect -1328 9210 -1288 13340
rect -968 9210 -928 13340
rect -1328 9170 -928 9210
rect -609 13340 -209 13380
rect -609 9210 -569 13340
rect -249 9210 -209 13340
rect -609 9170 -209 9210
rect 110 13340 510 13380
rect 110 9210 150 13340
rect 470 9210 510 13340
rect 110 9170 510 9210
rect 829 13340 1229 13380
rect 829 9210 869 13340
rect 1189 9210 1229 13340
rect 829 9170 1229 9210
rect 1548 13340 1948 13380
rect 1548 9210 1588 13340
rect 1908 9210 1948 13340
rect 1548 9170 1948 9210
rect 2267 13340 2667 13380
rect 2267 9210 2307 13340
rect 2627 9210 2667 13340
rect 2267 9170 2667 9210
rect -2766 8830 -2366 8870
rect -2766 4700 -2726 8830
rect -2406 4700 -2366 8830
rect -2766 4660 -2366 4700
rect -2047 8830 -1647 8870
rect -2047 4700 -2007 8830
rect -1687 4700 -1647 8830
rect -2047 4660 -1647 4700
rect -1328 8830 -928 8870
rect -1328 4700 -1288 8830
rect -968 4700 -928 8830
rect -1328 4660 -928 4700
rect -609 8830 -209 8870
rect -609 4700 -569 8830
rect -249 4700 -209 8830
rect -609 4660 -209 4700
rect 110 8830 510 8870
rect 110 4700 150 8830
rect 470 4700 510 8830
rect 110 4660 510 4700
rect 829 8830 1229 8870
rect 829 4700 869 8830
rect 1189 4700 1229 8830
rect 829 4660 1229 4700
rect 1548 8830 1948 8870
rect 1548 4700 1588 8830
rect 1908 4700 1948 8830
rect 1548 4660 1948 4700
rect 2267 8830 2667 8870
rect 2267 4700 2307 8830
rect 2627 4700 2667 8830
rect 2267 4660 2667 4700
rect -2766 4320 -2366 4360
rect -2766 190 -2726 4320
rect -2406 190 -2366 4320
rect -2766 150 -2366 190
rect -2047 4320 -1647 4360
rect -2047 190 -2007 4320
rect -1687 190 -1647 4320
rect -2047 150 -1647 190
rect -1328 4320 -928 4360
rect -1328 190 -1288 4320
rect -968 190 -928 4320
rect -1328 150 -928 190
rect -609 4320 -209 4360
rect -609 190 -569 4320
rect -249 190 -209 4320
rect -609 150 -209 190
rect 110 4320 510 4360
rect 110 190 150 4320
rect 470 190 510 4320
rect 110 150 510 190
rect 829 4320 1229 4360
rect 829 190 869 4320
rect 1189 190 1229 4320
rect 829 150 1229 190
rect 1548 4320 1948 4360
rect 1548 190 1588 4320
rect 1908 190 1948 4320
rect 1548 150 1948 190
rect 2267 4320 2667 4360
rect 2267 190 2307 4320
rect 2627 190 2667 4320
rect 2267 150 2667 190
rect -2766 -190 -2366 -150
rect -2766 -4320 -2726 -190
rect -2406 -4320 -2366 -190
rect -2766 -4360 -2366 -4320
rect -2047 -190 -1647 -150
rect -2047 -4320 -2007 -190
rect -1687 -4320 -1647 -190
rect -2047 -4360 -1647 -4320
rect -1328 -190 -928 -150
rect -1328 -4320 -1288 -190
rect -968 -4320 -928 -190
rect -1328 -4360 -928 -4320
rect -609 -190 -209 -150
rect -609 -4320 -569 -190
rect -249 -4320 -209 -190
rect -609 -4360 -209 -4320
rect 110 -190 510 -150
rect 110 -4320 150 -190
rect 470 -4320 510 -190
rect 110 -4360 510 -4320
rect 829 -190 1229 -150
rect 829 -4320 869 -190
rect 1189 -4320 1229 -190
rect 829 -4360 1229 -4320
rect 1548 -190 1948 -150
rect 1548 -4320 1588 -190
rect 1908 -4320 1948 -190
rect 1548 -4360 1948 -4320
rect 2267 -190 2667 -150
rect 2267 -4320 2307 -190
rect 2627 -4320 2667 -190
rect 2267 -4360 2667 -4320
rect -2766 -4700 -2366 -4660
rect -2766 -8830 -2726 -4700
rect -2406 -8830 -2366 -4700
rect -2766 -8870 -2366 -8830
rect -2047 -4700 -1647 -4660
rect -2047 -8830 -2007 -4700
rect -1687 -8830 -1647 -4700
rect -2047 -8870 -1647 -8830
rect -1328 -4700 -928 -4660
rect -1328 -8830 -1288 -4700
rect -968 -8830 -928 -4700
rect -1328 -8870 -928 -8830
rect -609 -4700 -209 -4660
rect -609 -8830 -569 -4700
rect -249 -8830 -209 -4700
rect -609 -8870 -209 -8830
rect 110 -4700 510 -4660
rect 110 -8830 150 -4700
rect 470 -8830 510 -4700
rect 110 -8870 510 -8830
rect 829 -4700 1229 -4660
rect 829 -8830 869 -4700
rect 1189 -8830 1229 -4700
rect 829 -8870 1229 -8830
rect 1548 -4700 1948 -4660
rect 1548 -8830 1588 -4700
rect 1908 -8830 1948 -4700
rect 1548 -8870 1948 -8830
rect 2267 -4700 2667 -4660
rect 2267 -8830 2307 -4700
rect 2627 -8830 2667 -4700
rect 2267 -8870 2667 -8830
rect -2766 -9210 -2366 -9170
rect -2766 -13340 -2726 -9210
rect -2406 -13340 -2366 -9210
rect -2766 -13380 -2366 -13340
rect -2047 -9210 -1647 -9170
rect -2047 -13340 -2007 -9210
rect -1687 -13340 -1647 -9210
rect -2047 -13380 -1647 -13340
rect -1328 -9210 -928 -9170
rect -1328 -13340 -1288 -9210
rect -968 -13340 -928 -9210
rect -1328 -13380 -928 -13340
rect -609 -9210 -209 -9170
rect -609 -13340 -569 -9210
rect -249 -13340 -209 -9210
rect -609 -13380 -209 -13340
rect 110 -9210 510 -9170
rect 110 -13340 150 -9210
rect 470 -13340 510 -9210
rect 110 -13380 510 -13340
rect 829 -9210 1229 -9170
rect 829 -13340 869 -9210
rect 1189 -13340 1229 -9210
rect 829 -13380 1229 -13340
rect 1548 -9210 1948 -9170
rect 1548 -13340 1588 -9210
rect 1908 -13340 1948 -9210
rect 1548 -13380 1948 -13340
rect 2267 -9210 2667 -9170
rect 2267 -13340 2307 -9210
rect 2627 -13340 2667 -9210
rect 2267 -13380 2667 -13340
rect -2766 -13720 -2366 -13680
rect -2766 -17850 -2726 -13720
rect -2406 -17850 -2366 -13720
rect -2766 -17890 -2366 -17850
rect -2047 -13720 -1647 -13680
rect -2047 -17850 -2007 -13720
rect -1687 -17850 -1647 -13720
rect -2047 -17890 -1647 -17850
rect -1328 -13720 -928 -13680
rect -1328 -17850 -1288 -13720
rect -968 -17850 -928 -13720
rect -1328 -17890 -928 -17850
rect -609 -13720 -209 -13680
rect -609 -17850 -569 -13720
rect -249 -17850 -209 -13720
rect -609 -17890 -209 -17850
rect 110 -13720 510 -13680
rect 110 -17850 150 -13720
rect 470 -17850 510 -13720
rect 110 -17890 510 -17850
rect 829 -13720 1229 -13680
rect 829 -17850 869 -13720
rect 1189 -17850 1229 -13720
rect 829 -17890 1229 -17850
rect 1548 -13720 1948 -13680
rect 1548 -17850 1588 -13720
rect 1908 -17850 1948 -13720
rect 1548 -17890 1948 -17850
rect 2267 -13720 2667 -13680
rect 2267 -17850 2307 -13720
rect 2627 -17850 2667 -13720
rect 2267 -17890 2667 -17850
rect -2766 -18230 -2366 -18190
rect -2766 -22360 -2726 -18230
rect -2406 -22360 -2366 -18230
rect -2766 -22400 -2366 -22360
rect -2047 -18230 -1647 -18190
rect -2047 -22360 -2007 -18230
rect -1687 -22360 -1647 -18230
rect -2047 -22400 -1647 -22360
rect -1328 -18230 -928 -18190
rect -1328 -22360 -1288 -18230
rect -968 -22360 -928 -18230
rect -1328 -22400 -928 -22360
rect -609 -18230 -209 -18190
rect -609 -22360 -569 -18230
rect -249 -22360 -209 -18230
rect -609 -22400 -209 -22360
rect 110 -18230 510 -18190
rect 110 -22360 150 -18230
rect 470 -22360 510 -18230
rect 110 -22400 510 -22360
rect 829 -18230 1229 -18190
rect 829 -22360 869 -18230
rect 1189 -22360 1229 -18230
rect 829 -22400 1229 -22360
rect 1548 -18230 1948 -18190
rect 1548 -22360 1588 -18230
rect 1908 -22360 1948 -18230
rect 1548 -22400 1948 -22360
rect 2267 -18230 2667 -18190
rect 2267 -22360 2307 -18230
rect 2627 -22360 2667 -18230
rect 2267 -22400 2667 -22360
rect -2766 -22740 -2366 -22700
rect -2766 -26870 -2726 -22740
rect -2406 -26870 -2366 -22740
rect -2766 -26910 -2366 -26870
rect -2047 -22740 -1647 -22700
rect -2047 -26870 -2007 -22740
rect -1687 -26870 -1647 -22740
rect -2047 -26910 -1647 -26870
rect -1328 -22740 -928 -22700
rect -1328 -26870 -1288 -22740
rect -968 -26870 -928 -22740
rect -1328 -26910 -928 -26870
rect -609 -22740 -209 -22700
rect -609 -26870 -569 -22740
rect -249 -26870 -209 -22740
rect -609 -26910 -209 -26870
rect 110 -22740 510 -22700
rect 110 -26870 150 -22740
rect 470 -26870 510 -22740
rect 110 -26910 510 -26870
rect 829 -22740 1229 -22700
rect 829 -26870 869 -22740
rect 1189 -26870 1229 -22740
rect 829 -26910 1229 -26870
rect 1548 -22740 1948 -22700
rect 1548 -26870 1588 -22740
rect 1908 -26870 1948 -22740
rect 1548 -26910 1948 -26870
rect 2267 -22740 2667 -22700
rect 2267 -26870 2307 -22740
rect 2627 -26870 2667 -22740
rect 2267 -26910 2667 -26870
rect -2766 -27250 -2366 -27210
rect -2766 -31380 -2726 -27250
rect -2406 -31380 -2366 -27250
rect -2766 -31420 -2366 -31380
rect -2047 -27250 -1647 -27210
rect -2047 -31380 -2007 -27250
rect -1687 -31380 -1647 -27250
rect -2047 -31420 -1647 -31380
rect -1328 -27250 -928 -27210
rect -1328 -31380 -1288 -27250
rect -968 -31380 -928 -27250
rect -1328 -31420 -928 -31380
rect -609 -27250 -209 -27210
rect -609 -31380 -569 -27250
rect -249 -31380 -209 -27250
rect -609 -31420 -209 -31380
rect 110 -27250 510 -27210
rect 110 -31380 150 -27250
rect 470 -31380 510 -27250
rect 110 -31420 510 -31380
rect 829 -27250 1229 -27210
rect 829 -31380 869 -27250
rect 1189 -31380 1229 -27250
rect 829 -31420 1229 -31380
rect 1548 -27250 1948 -27210
rect 1548 -31380 1588 -27250
rect 1908 -31380 1948 -27250
rect 1548 -31420 1948 -31380
rect 2267 -27250 2667 -27210
rect 2267 -31380 2307 -27250
rect 2627 -31380 2667 -27250
rect 2267 -31420 2667 -31380
rect -2766 -31760 -2366 -31720
rect -2766 -35890 -2726 -31760
rect -2406 -35890 -2366 -31760
rect -2766 -35930 -2366 -35890
rect -2047 -31760 -1647 -31720
rect -2047 -35890 -2007 -31760
rect -1687 -35890 -1647 -31760
rect -2047 -35930 -1647 -35890
rect -1328 -31760 -928 -31720
rect -1328 -35890 -1288 -31760
rect -968 -35890 -928 -31760
rect -1328 -35930 -928 -35890
rect -609 -31760 -209 -31720
rect -609 -35890 -569 -31760
rect -249 -35890 -209 -31760
rect -609 -35930 -209 -35890
rect 110 -31760 510 -31720
rect 110 -35890 150 -31760
rect 470 -35890 510 -31760
rect 110 -35930 510 -35890
rect 829 -31760 1229 -31720
rect 829 -35890 869 -31760
rect 1189 -35890 1229 -31760
rect 829 -35930 1229 -35890
rect 1548 -31760 1948 -31720
rect 1548 -35890 1588 -31760
rect 1908 -35890 1948 -31760
rect 1548 -35930 1948 -35890
rect 2267 -31760 2667 -31720
rect 2267 -35890 2307 -31760
rect 2627 -35890 2667 -31760
rect 2267 -35930 2667 -35890
<< mimcapcontact >>
rect -2726 31760 -2406 35890
rect -2007 31760 -1687 35890
rect -1288 31760 -968 35890
rect -569 31760 -249 35890
rect 150 31760 470 35890
rect 869 31760 1189 35890
rect 1588 31760 1908 35890
rect 2307 31760 2627 35890
rect -2726 27250 -2406 31380
rect -2007 27250 -1687 31380
rect -1288 27250 -968 31380
rect -569 27250 -249 31380
rect 150 27250 470 31380
rect 869 27250 1189 31380
rect 1588 27250 1908 31380
rect 2307 27250 2627 31380
rect -2726 22740 -2406 26870
rect -2007 22740 -1687 26870
rect -1288 22740 -968 26870
rect -569 22740 -249 26870
rect 150 22740 470 26870
rect 869 22740 1189 26870
rect 1588 22740 1908 26870
rect 2307 22740 2627 26870
rect -2726 18230 -2406 22360
rect -2007 18230 -1687 22360
rect -1288 18230 -968 22360
rect -569 18230 -249 22360
rect 150 18230 470 22360
rect 869 18230 1189 22360
rect 1588 18230 1908 22360
rect 2307 18230 2627 22360
rect -2726 13720 -2406 17850
rect -2007 13720 -1687 17850
rect -1288 13720 -968 17850
rect -569 13720 -249 17850
rect 150 13720 470 17850
rect 869 13720 1189 17850
rect 1588 13720 1908 17850
rect 2307 13720 2627 17850
rect -2726 9210 -2406 13340
rect -2007 9210 -1687 13340
rect -1288 9210 -968 13340
rect -569 9210 -249 13340
rect 150 9210 470 13340
rect 869 9210 1189 13340
rect 1588 9210 1908 13340
rect 2307 9210 2627 13340
rect -2726 4700 -2406 8830
rect -2007 4700 -1687 8830
rect -1288 4700 -968 8830
rect -569 4700 -249 8830
rect 150 4700 470 8830
rect 869 4700 1189 8830
rect 1588 4700 1908 8830
rect 2307 4700 2627 8830
rect -2726 190 -2406 4320
rect -2007 190 -1687 4320
rect -1288 190 -968 4320
rect -569 190 -249 4320
rect 150 190 470 4320
rect 869 190 1189 4320
rect 1588 190 1908 4320
rect 2307 190 2627 4320
rect -2726 -4320 -2406 -190
rect -2007 -4320 -1687 -190
rect -1288 -4320 -968 -190
rect -569 -4320 -249 -190
rect 150 -4320 470 -190
rect 869 -4320 1189 -190
rect 1588 -4320 1908 -190
rect 2307 -4320 2627 -190
rect -2726 -8830 -2406 -4700
rect -2007 -8830 -1687 -4700
rect -1288 -8830 -968 -4700
rect -569 -8830 -249 -4700
rect 150 -8830 470 -4700
rect 869 -8830 1189 -4700
rect 1588 -8830 1908 -4700
rect 2307 -8830 2627 -4700
rect -2726 -13340 -2406 -9210
rect -2007 -13340 -1687 -9210
rect -1288 -13340 -968 -9210
rect -569 -13340 -249 -9210
rect 150 -13340 470 -9210
rect 869 -13340 1189 -9210
rect 1588 -13340 1908 -9210
rect 2307 -13340 2627 -9210
rect -2726 -17850 -2406 -13720
rect -2007 -17850 -1687 -13720
rect -1288 -17850 -968 -13720
rect -569 -17850 -249 -13720
rect 150 -17850 470 -13720
rect 869 -17850 1189 -13720
rect 1588 -17850 1908 -13720
rect 2307 -17850 2627 -13720
rect -2726 -22360 -2406 -18230
rect -2007 -22360 -1687 -18230
rect -1288 -22360 -968 -18230
rect -569 -22360 -249 -18230
rect 150 -22360 470 -18230
rect 869 -22360 1189 -18230
rect 1588 -22360 1908 -18230
rect 2307 -22360 2627 -18230
rect -2726 -26870 -2406 -22740
rect -2007 -26870 -1687 -22740
rect -1288 -26870 -968 -22740
rect -569 -26870 -249 -22740
rect 150 -26870 470 -22740
rect 869 -26870 1189 -22740
rect 1588 -26870 1908 -22740
rect 2307 -26870 2627 -22740
rect -2726 -31380 -2406 -27250
rect -2007 -31380 -1687 -27250
rect -1288 -31380 -968 -27250
rect -569 -31380 -249 -27250
rect 150 -31380 470 -27250
rect 869 -31380 1189 -27250
rect 1588 -31380 1908 -27250
rect 2307 -31380 2627 -27250
rect -2726 -35890 -2406 -31760
rect -2007 -35890 -1687 -31760
rect -1288 -35890 -968 -31760
rect -569 -35890 -249 -31760
rect 150 -35890 470 -31760
rect 869 -35890 1189 -31760
rect 1588 -35890 1908 -31760
rect 2307 -35890 2627 -31760
<< metal4 >>
rect -2618 35891 -2514 36080
rect -2298 36018 -2194 36080
rect -2298 36002 -2171 36018
rect -2727 35890 -2405 35891
rect -2727 31760 -2726 35890
rect -2406 31760 -2405 35890
rect -2727 31759 -2405 31760
rect -2618 31381 -2514 31759
rect -2298 31648 -2251 36002
rect -2187 31648 -2171 36002
rect -1899 35891 -1795 36080
rect -1579 36018 -1475 36080
rect -1579 36002 -1452 36018
rect -2008 35890 -1686 35891
rect -2008 31760 -2007 35890
rect -1687 31760 -1686 35890
rect -2008 31759 -1686 31760
rect -2298 31632 -2171 31648
rect -2298 31508 -2194 31632
rect -2298 31492 -2171 31508
rect -2727 31380 -2405 31381
rect -2727 27250 -2726 31380
rect -2406 27250 -2405 31380
rect -2727 27249 -2405 27250
rect -2618 26871 -2514 27249
rect -2298 27138 -2251 31492
rect -2187 27138 -2171 31492
rect -1899 31381 -1795 31759
rect -1579 31648 -1532 36002
rect -1468 31648 -1452 36002
rect -1180 35891 -1076 36080
rect -860 36018 -756 36080
rect -860 36002 -733 36018
rect -1289 35890 -967 35891
rect -1289 31760 -1288 35890
rect -968 31760 -967 35890
rect -1289 31759 -967 31760
rect -1579 31632 -1452 31648
rect -1579 31508 -1475 31632
rect -1579 31492 -1452 31508
rect -2008 31380 -1686 31381
rect -2008 27250 -2007 31380
rect -1687 27250 -1686 31380
rect -2008 27249 -1686 27250
rect -2298 27122 -2171 27138
rect -2298 26998 -2194 27122
rect -2298 26982 -2171 26998
rect -2727 26870 -2405 26871
rect -2727 22740 -2726 26870
rect -2406 22740 -2405 26870
rect -2727 22739 -2405 22740
rect -2618 22361 -2514 22739
rect -2298 22628 -2251 26982
rect -2187 22628 -2171 26982
rect -1899 26871 -1795 27249
rect -1579 27138 -1532 31492
rect -1468 27138 -1452 31492
rect -1180 31381 -1076 31759
rect -860 31648 -813 36002
rect -749 31648 -733 36002
rect -461 35891 -357 36080
rect -141 36018 -37 36080
rect -141 36002 -14 36018
rect -570 35890 -248 35891
rect -570 31760 -569 35890
rect -249 31760 -248 35890
rect -570 31759 -248 31760
rect -860 31632 -733 31648
rect -860 31508 -756 31632
rect -860 31492 -733 31508
rect -1289 31380 -967 31381
rect -1289 27250 -1288 31380
rect -968 27250 -967 31380
rect -1289 27249 -967 27250
rect -1579 27122 -1452 27138
rect -1579 26998 -1475 27122
rect -1579 26982 -1452 26998
rect -2008 26870 -1686 26871
rect -2008 22740 -2007 26870
rect -1687 22740 -1686 26870
rect -2008 22739 -1686 22740
rect -2298 22612 -2171 22628
rect -2298 22488 -2194 22612
rect -2298 22472 -2171 22488
rect -2727 22360 -2405 22361
rect -2727 18230 -2726 22360
rect -2406 18230 -2405 22360
rect -2727 18229 -2405 18230
rect -2618 17851 -2514 18229
rect -2298 18118 -2251 22472
rect -2187 18118 -2171 22472
rect -1899 22361 -1795 22739
rect -1579 22628 -1532 26982
rect -1468 22628 -1452 26982
rect -1180 26871 -1076 27249
rect -860 27138 -813 31492
rect -749 27138 -733 31492
rect -461 31381 -357 31759
rect -141 31648 -94 36002
rect -30 31648 -14 36002
rect 258 35891 362 36080
rect 578 36018 682 36080
rect 578 36002 705 36018
rect 149 35890 471 35891
rect 149 31760 150 35890
rect 470 31760 471 35890
rect 149 31759 471 31760
rect -141 31632 -14 31648
rect -141 31508 -37 31632
rect -141 31492 -14 31508
rect -570 31380 -248 31381
rect -570 27250 -569 31380
rect -249 27250 -248 31380
rect -570 27249 -248 27250
rect -860 27122 -733 27138
rect -860 26998 -756 27122
rect -860 26982 -733 26998
rect -1289 26870 -967 26871
rect -1289 22740 -1288 26870
rect -968 22740 -967 26870
rect -1289 22739 -967 22740
rect -1579 22612 -1452 22628
rect -1579 22488 -1475 22612
rect -1579 22472 -1452 22488
rect -2008 22360 -1686 22361
rect -2008 18230 -2007 22360
rect -1687 18230 -1686 22360
rect -2008 18229 -1686 18230
rect -2298 18102 -2171 18118
rect -2298 17978 -2194 18102
rect -2298 17962 -2171 17978
rect -2727 17850 -2405 17851
rect -2727 13720 -2726 17850
rect -2406 13720 -2405 17850
rect -2727 13719 -2405 13720
rect -2618 13341 -2514 13719
rect -2298 13608 -2251 17962
rect -2187 13608 -2171 17962
rect -1899 17851 -1795 18229
rect -1579 18118 -1532 22472
rect -1468 18118 -1452 22472
rect -1180 22361 -1076 22739
rect -860 22628 -813 26982
rect -749 22628 -733 26982
rect -461 26871 -357 27249
rect -141 27138 -94 31492
rect -30 27138 -14 31492
rect 258 31381 362 31759
rect 578 31648 625 36002
rect 689 31648 705 36002
rect 977 35891 1081 36080
rect 1297 36018 1401 36080
rect 1297 36002 1424 36018
rect 868 35890 1190 35891
rect 868 31760 869 35890
rect 1189 31760 1190 35890
rect 868 31759 1190 31760
rect 578 31632 705 31648
rect 578 31508 682 31632
rect 578 31492 705 31508
rect 149 31380 471 31381
rect 149 27250 150 31380
rect 470 27250 471 31380
rect 149 27249 471 27250
rect -141 27122 -14 27138
rect -141 26998 -37 27122
rect -141 26982 -14 26998
rect -570 26870 -248 26871
rect -570 22740 -569 26870
rect -249 22740 -248 26870
rect -570 22739 -248 22740
rect -860 22612 -733 22628
rect -860 22488 -756 22612
rect -860 22472 -733 22488
rect -1289 22360 -967 22361
rect -1289 18230 -1288 22360
rect -968 18230 -967 22360
rect -1289 18229 -967 18230
rect -1579 18102 -1452 18118
rect -1579 17978 -1475 18102
rect -1579 17962 -1452 17978
rect -2008 17850 -1686 17851
rect -2008 13720 -2007 17850
rect -1687 13720 -1686 17850
rect -2008 13719 -1686 13720
rect -2298 13592 -2171 13608
rect -2298 13468 -2194 13592
rect -2298 13452 -2171 13468
rect -2727 13340 -2405 13341
rect -2727 9210 -2726 13340
rect -2406 9210 -2405 13340
rect -2727 9209 -2405 9210
rect -2618 8831 -2514 9209
rect -2298 9098 -2251 13452
rect -2187 9098 -2171 13452
rect -1899 13341 -1795 13719
rect -1579 13608 -1532 17962
rect -1468 13608 -1452 17962
rect -1180 17851 -1076 18229
rect -860 18118 -813 22472
rect -749 18118 -733 22472
rect -461 22361 -357 22739
rect -141 22628 -94 26982
rect -30 22628 -14 26982
rect 258 26871 362 27249
rect 578 27138 625 31492
rect 689 27138 705 31492
rect 977 31381 1081 31759
rect 1297 31648 1344 36002
rect 1408 31648 1424 36002
rect 1696 35891 1800 36080
rect 2016 36018 2120 36080
rect 2016 36002 2143 36018
rect 1587 35890 1909 35891
rect 1587 31760 1588 35890
rect 1908 31760 1909 35890
rect 1587 31759 1909 31760
rect 1297 31632 1424 31648
rect 1297 31508 1401 31632
rect 1297 31492 1424 31508
rect 868 31380 1190 31381
rect 868 27250 869 31380
rect 1189 27250 1190 31380
rect 868 27249 1190 27250
rect 578 27122 705 27138
rect 578 26998 682 27122
rect 578 26982 705 26998
rect 149 26870 471 26871
rect 149 22740 150 26870
rect 470 22740 471 26870
rect 149 22739 471 22740
rect -141 22612 -14 22628
rect -141 22488 -37 22612
rect -141 22472 -14 22488
rect -570 22360 -248 22361
rect -570 18230 -569 22360
rect -249 18230 -248 22360
rect -570 18229 -248 18230
rect -860 18102 -733 18118
rect -860 17978 -756 18102
rect -860 17962 -733 17978
rect -1289 17850 -967 17851
rect -1289 13720 -1288 17850
rect -968 13720 -967 17850
rect -1289 13719 -967 13720
rect -1579 13592 -1452 13608
rect -1579 13468 -1475 13592
rect -1579 13452 -1452 13468
rect -2008 13340 -1686 13341
rect -2008 9210 -2007 13340
rect -1687 9210 -1686 13340
rect -2008 9209 -1686 9210
rect -2298 9082 -2171 9098
rect -2298 8958 -2194 9082
rect -2298 8942 -2171 8958
rect -2727 8830 -2405 8831
rect -2727 4700 -2726 8830
rect -2406 4700 -2405 8830
rect -2727 4699 -2405 4700
rect -2618 4321 -2514 4699
rect -2298 4588 -2251 8942
rect -2187 4588 -2171 8942
rect -1899 8831 -1795 9209
rect -1579 9098 -1532 13452
rect -1468 9098 -1452 13452
rect -1180 13341 -1076 13719
rect -860 13608 -813 17962
rect -749 13608 -733 17962
rect -461 17851 -357 18229
rect -141 18118 -94 22472
rect -30 18118 -14 22472
rect 258 22361 362 22739
rect 578 22628 625 26982
rect 689 22628 705 26982
rect 977 26871 1081 27249
rect 1297 27138 1344 31492
rect 1408 27138 1424 31492
rect 1696 31381 1800 31759
rect 2016 31648 2063 36002
rect 2127 31648 2143 36002
rect 2415 35891 2519 36080
rect 2735 36018 2839 36080
rect 2735 36002 2862 36018
rect 2306 35890 2628 35891
rect 2306 31760 2307 35890
rect 2627 31760 2628 35890
rect 2306 31759 2628 31760
rect 2016 31632 2143 31648
rect 2016 31508 2120 31632
rect 2016 31492 2143 31508
rect 1587 31380 1909 31381
rect 1587 27250 1588 31380
rect 1908 27250 1909 31380
rect 1587 27249 1909 27250
rect 1297 27122 1424 27138
rect 1297 26998 1401 27122
rect 1297 26982 1424 26998
rect 868 26870 1190 26871
rect 868 22740 869 26870
rect 1189 22740 1190 26870
rect 868 22739 1190 22740
rect 578 22612 705 22628
rect 578 22488 682 22612
rect 578 22472 705 22488
rect 149 22360 471 22361
rect 149 18230 150 22360
rect 470 18230 471 22360
rect 149 18229 471 18230
rect -141 18102 -14 18118
rect -141 17978 -37 18102
rect -141 17962 -14 17978
rect -570 17850 -248 17851
rect -570 13720 -569 17850
rect -249 13720 -248 17850
rect -570 13719 -248 13720
rect -860 13592 -733 13608
rect -860 13468 -756 13592
rect -860 13452 -733 13468
rect -1289 13340 -967 13341
rect -1289 9210 -1288 13340
rect -968 9210 -967 13340
rect -1289 9209 -967 9210
rect -1579 9082 -1452 9098
rect -1579 8958 -1475 9082
rect -1579 8942 -1452 8958
rect -2008 8830 -1686 8831
rect -2008 4700 -2007 8830
rect -1687 4700 -1686 8830
rect -2008 4699 -1686 4700
rect -2298 4572 -2171 4588
rect -2298 4448 -2194 4572
rect -2298 4432 -2171 4448
rect -2727 4320 -2405 4321
rect -2727 190 -2726 4320
rect -2406 190 -2405 4320
rect -2727 189 -2405 190
rect -2618 -189 -2514 189
rect -2298 78 -2251 4432
rect -2187 78 -2171 4432
rect -1899 4321 -1795 4699
rect -1579 4588 -1532 8942
rect -1468 4588 -1452 8942
rect -1180 8831 -1076 9209
rect -860 9098 -813 13452
rect -749 9098 -733 13452
rect -461 13341 -357 13719
rect -141 13608 -94 17962
rect -30 13608 -14 17962
rect 258 17851 362 18229
rect 578 18118 625 22472
rect 689 18118 705 22472
rect 977 22361 1081 22739
rect 1297 22628 1344 26982
rect 1408 22628 1424 26982
rect 1696 26871 1800 27249
rect 2016 27138 2063 31492
rect 2127 27138 2143 31492
rect 2415 31381 2519 31759
rect 2735 31648 2782 36002
rect 2846 31648 2862 36002
rect 2735 31632 2862 31648
rect 2735 31508 2839 31632
rect 2735 31492 2862 31508
rect 2306 31380 2628 31381
rect 2306 27250 2307 31380
rect 2627 27250 2628 31380
rect 2306 27249 2628 27250
rect 2016 27122 2143 27138
rect 2016 26998 2120 27122
rect 2016 26982 2143 26998
rect 1587 26870 1909 26871
rect 1587 22740 1588 26870
rect 1908 22740 1909 26870
rect 1587 22739 1909 22740
rect 1297 22612 1424 22628
rect 1297 22488 1401 22612
rect 1297 22472 1424 22488
rect 868 22360 1190 22361
rect 868 18230 869 22360
rect 1189 18230 1190 22360
rect 868 18229 1190 18230
rect 578 18102 705 18118
rect 578 17978 682 18102
rect 578 17962 705 17978
rect 149 17850 471 17851
rect 149 13720 150 17850
rect 470 13720 471 17850
rect 149 13719 471 13720
rect -141 13592 -14 13608
rect -141 13468 -37 13592
rect -141 13452 -14 13468
rect -570 13340 -248 13341
rect -570 9210 -569 13340
rect -249 9210 -248 13340
rect -570 9209 -248 9210
rect -860 9082 -733 9098
rect -860 8958 -756 9082
rect -860 8942 -733 8958
rect -1289 8830 -967 8831
rect -1289 4700 -1288 8830
rect -968 4700 -967 8830
rect -1289 4699 -967 4700
rect -1579 4572 -1452 4588
rect -1579 4448 -1475 4572
rect -1579 4432 -1452 4448
rect -2008 4320 -1686 4321
rect -2008 190 -2007 4320
rect -1687 190 -1686 4320
rect -2008 189 -1686 190
rect -2298 62 -2171 78
rect -2298 -62 -2194 62
rect -2298 -78 -2171 -62
rect -2727 -190 -2405 -189
rect -2727 -4320 -2726 -190
rect -2406 -4320 -2405 -190
rect -2727 -4321 -2405 -4320
rect -2618 -4699 -2514 -4321
rect -2298 -4432 -2251 -78
rect -2187 -4432 -2171 -78
rect -1899 -189 -1795 189
rect -1579 78 -1532 4432
rect -1468 78 -1452 4432
rect -1180 4321 -1076 4699
rect -860 4588 -813 8942
rect -749 4588 -733 8942
rect -461 8831 -357 9209
rect -141 9098 -94 13452
rect -30 9098 -14 13452
rect 258 13341 362 13719
rect 578 13608 625 17962
rect 689 13608 705 17962
rect 977 17851 1081 18229
rect 1297 18118 1344 22472
rect 1408 18118 1424 22472
rect 1696 22361 1800 22739
rect 2016 22628 2063 26982
rect 2127 22628 2143 26982
rect 2415 26871 2519 27249
rect 2735 27138 2782 31492
rect 2846 27138 2862 31492
rect 2735 27122 2862 27138
rect 2735 26998 2839 27122
rect 2735 26982 2862 26998
rect 2306 26870 2628 26871
rect 2306 22740 2307 26870
rect 2627 22740 2628 26870
rect 2306 22739 2628 22740
rect 2016 22612 2143 22628
rect 2016 22488 2120 22612
rect 2016 22472 2143 22488
rect 1587 22360 1909 22361
rect 1587 18230 1588 22360
rect 1908 18230 1909 22360
rect 1587 18229 1909 18230
rect 1297 18102 1424 18118
rect 1297 17978 1401 18102
rect 1297 17962 1424 17978
rect 868 17850 1190 17851
rect 868 13720 869 17850
rect 1189 13720 1190 17850
rect 868 13719 1190 13720
rect 578 13592 705 13608
rect 578 13468 682 13592
rect 578 13452 705 13468
rect 149 13340 471 13341
rect 149 9210 150 13340
rect 470 9210 471 13340
rect 149 9209 471 9210
rect -141 9082 -14 9098
rect -141 8958 -37 9082
rect -141 8942 -14 8958
rect -570 8830 -248 8831
rect -570 4700 -569 8830
rect -249 4700 -248 8830
rect -570 4699 -248 4700
rect -860 4572 -733 4588
rect -860 4448 -756 4572
rect -860 4432 -733 4448
rect -1289 4320 -967 4321
rect -1289 190 -1288 4320
rect -968 190 -967 4320
rect -1289 189 -967 190
rect -1579 62 -1452 78
rect -1579 -62 -1475 62
rect -1579 -78 -1452 -62
rect -2008 -190 -1686 -189
rect -2008 -4320 -2007 -190
rect -1687 -4320 -1686 -190
rect -2008 -4321 -1686 -4320
rect -2298 -4448 -2171 -4432
rect -2298 -4572 -2194 -4448
rect -2298 -4588 -2171 -4572
rect -2727 -4700 -2405 -4699
rect -2727 -8830 -2726 -4700
rect -2406 -8830 -2405 -4700
rect -2727 -8831 -2405 -8830
rect -2618 -9209 -2514 -8831
rect -2298 -8942 -2251 -4588
rect -2187 -8942 -2171 -4588
rect -1899 -4699 -1795 -4321
rect -1579 -4432 -1532 -78
rect -1468 -4432 -1452 -78
rect -1180 -189 -1076 189
rect -860 78 -813 4432
rect -749 78 -733 4432
rect -461 4321 -357 4699
rect -141 4588 -94 8942
rect -30 4588 -14 8942
rect 258 8831 362 9209
rect 578 9098 625 13452
rect 689 9098 705 13452
rect 977 13341 1081 13719
rect 1297 13608 1344 17962
rect 1408 13608 1424 17962
rect 1696 17851 1800 18229
rect 2016 18118 2063 22472
rect 2127 18118 2143 22472
rect 2415 22361 2519 22739
rect 2735 22628 2782 26982
rect 2846 22628 2862 26982
rect 2735 22612 2862 22628
rect 2735 22488 2839 22612
rect 2735 22472 2862 22488
rect 2306 22360 2628 22361
rect 2306 18230 2307 22360
rect 2627 18230 2628 22360
rect 2306 18229 2628 18230
rect 2016 18102 2143 18118
rect 2016 17978 2120 18102
rect 2016 17962 2143 17978
rect 1587 17850 1909 17851
rect 1587 13720 1588 17850
rect 1908 13720 1909 17850
rect 1587 13719 1909 13720
rect 1297 13592 1424 13608
rect 1297 13468 1401 13592
rect 1297 13452 1424 13468
rect 868 13340 1190 13341
rect 868 9210 869 13340
rect 1189 9210 1190 13340
rect 868 9209 1190 9210
rect 578 9082 705 9098
rect 578 8958 682 9082
rect 578 8942 705 8958
rect 149 8830 471 8831
rect 149 4700 150 8830
rect 470 4700 471 8830
rect 149 4699 471 4700
rect -141 4572 -14 4588
rect -141 4448 -37 4572
rect -141 4432 -14 4448
rect -570 4320 -248 4321
rect -570 190 -569 4320
rect -249 190 -248 4320
rect -570 189 -248 190
rect -860 62 -733 78
rect -860 -62 -756 62
rect -860 -78 -733 -62
rect -1289 -190 -967 -189
rect -1289 -4320 -1288 -190
rect -968 -4320 -967 -190
rect -1289 -4321 -967 -4320
rect -1579 -4448 -1452 -4432
rect -1579 -4572 -1475 -4448
rect -1579 -4588 -1452 -4572
rect -2008 -4700 -1686 -4699
rect -2008 -8830 -2007 -4700
rect -1687 -8830 -1686 -4700
rect -2008 -8831 -1686 -8830
rect -2298 -8958 -2171 -8942
rect -2298 -9082 -2194 -8958
rect -2298 -9098 -2171 -9082
rect -2727 -9210 -2405 -9209
rect -2727 -13340 -2726 -9210
rect -2406 -13340 -2405 -9210
rect -2727 -13341 -2405 -13340
rect -2618 -13719 -2514 -13341
rect -2298 -13452 -2251 -9098
rect -2187 -13452 -2171 -9098
rect -1899 -9209 -1795 -8831
rect -1579 -8942 -1532 -4588
rect -1468 -8942 -1452 -4588
rect -1180 -4699 -1076 -4321
rect -860 -4432 -813 -78
rect -749 -4432 -733 -78
rect -461 -189 -357 189
rect -141 78 -94 4432
rect -30 78 -14 4432
rect 258 4321 362 4699
rect 578 4588 625 8942
rect 689 4588 705 8942
rect 977 8831 1081 9209
rect 1297 9098 1344 13452
rect 1408 9098 1424 13452
rect 1696 13341 1800 13719
rect 2016 13608 2063 17962
rect 2127 13608 2143 17962
rect 2415 17851 2519 18229
rect 2735 18118 2782 22472
rect 2846 18118 2862 22472
rect 2735 18102 2862 18118
rect 2735 17978 2839 18102
rect 2735 17962 2862 17978
rect 2306 17850 2628 17851
rect 2306 13720 2307 17850
rect 2627 13720 2628 17850
rect 2306 13719 2628 13720
rect 2016 13592 2143 13608
rect 2016 13468 2120 13592
rect 2016 13452 2143 13468
rect 1587 13340 1909 13341
rect 1587 9210 1588 13340
rect 1908 9210 1909 13340
rect 1587 9209 1909 9210
rect 1297 9082 1424 9098
rect 1297 8958 1401 9082
rect 1297 8942 1424 8958
rect 868 8830 1190 8831
rect 868 4700 869 8830
rect 1189 4700 1190 8830
rect 868 4699 1190 4700
rect 578 4572 705 4588
rect 578 4448 682 4572
rect 578 4432 705 4448
rect 149 4320 471 4321
rect 149 190 150 4320
rect 470 190 471 4320
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -4320 -569 -190
rect -249 -4320 -248 -190
rect -570 -4321 -248 -4320
rect -860 -4448 -733 -4432
rect -860 -4572 -756 -4448
rect -860 -4588 -733 -4572
rect -1289 -4700 -967 -4699
rect -1289 -8830 -1288 -4700
rect -968 -8830 -967 -4700
rect -1289 -8831 -967 -8830
rect -1579 -8958 -1452 -8942
rect -1579 -9082 -1475 -8958
rect -1579 -9098 -1452 -9082
rect -2008 -9210 -1686 -9209
rect -2008 -13340 -2007 -9210
rect -1687 -13340 -1686 -9210
rect -2008 -13341 -1686 -13340
rect -2298 -13468 -2171 -13452
rect -2298 -13592 -2194 -13468
rect -2298 -13608 -2171 -13592
rect -2727 -13720 -2405 -13719
rect -2727 -17850 -2726 -13720
rect -2406 -17850 -2405 -13720
rect -2727 -17851 -2405 -17850
rect -2618 -18229 -2514 -17851
rect -2298 -17962 -2251 -13608
rect -2187 -17962 -2171 -13608
rect -1899 -13719 -1795 -13341
rect -1579 -13452 -1532 -9098
rect -1468 -13452 -1452 -9098
rect -1180 -9209 -1076 -8831
rect -860 -8942 -813 -4588
rect -749 -8942 -733 -4588
rect -461 -4699 -357 -4321
rect -141 -4432 -94 -78
rect -30 -4432 -14 -78
rect 258 -189 362 189
rect 578 78 625 4432
rect 689 78 705 4432
rect 977 4321 1081 4699
rect 1297 4588 1344 8942
rect 1408 4588 1424 8942
rect 1696 8831 1800 9209
rect 2016 9098 2063 13452
rect 2127 9098 2143 13452
rect 2415 13341 2519 13719
rect 2735 13608 2782 17962
rect 2846 13608 2862 17962
rect 2735 13592 2862 13608
rect 2735 13468 2839 13592
rect 2735 13452 2862 13468
rect 2306 13340 2628 13341
rect 2306 9210 2307 13340
rect 2627 9210 2628 13340
rect 2306 9209 2628 9210
rect 2016 9082 2143 9098
rect 2016 8958 2120 9082
rect 2016 8942 2143 8958
rect 1587 8830 1909 8831
rect 1587 4700 1588 8830
rect 1908 4700 1909 8830
rect 1587 4699 1909 4700
rect 1297 4572 1424 4588
rect 1297 4448 1401 4572
rect 1297 4432 1424 4448
rect 868 4320 1190 4321
rect 868 190 869 4320
rect 1189 190 1190 4320
rect 868 189 1190 190
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -4320 150 -190
rect 470 -4320 471 -190
rect 149 -4321 471 -4320
rect -141 -4448 -14 -4432
rect -141 -4572 -37 -4448
rect -141 -4588 -14 -4572
rect -570 -4700 -248 -4699
rect -570 -8830 -569 -4700
rect -249 -8830 -248 -4700
rect -570 -8831 -248 -8830
rect -860 -8958 -733 -8942
rect -860 -9082 -756 -8958
rect -860 -9098 -733 -9082
rect -1289 -9210 -967 -9209
rect -1289 -13340 -1288 -9210
rect -968 -13340 -967 -9210
rect -1289 -13341 -967 -13340
rect -1579 -13468 -1452 -13452
rect -1579 -13592 -1475 -13468
rect -1579 -13608 -1452 -13592
rect -2008 -13720 -1686 -13719
rect -2008 -17850 -2007 -13720
rect -1687 -17850 -1686 -13720
rect -2008 -17851 -1686 -17850
rect -2298 -17978 -2171 -17962
rect -2298 -18102 -2194 -17978
rect -2298 -18118 -2171 -18102
rect -2727 -18230 -2405 -18229
rect -2727 -22360 -2726 -18230
rect -2406 -22360 -2405 -18230
rect -2727 -22361 -2405 -22360
rect -2618 -22739 -2514 -22361
rect -2298 -22472 -2251 -18118
rect -2187 -22472 -2171 -18118
rect -1899 -18229 -1795 -17851
rect -1579 -17962 -1532 -13608
rect -1468 -17962 -1452 -13608
rect -1180 -13719 -1076 -13341
rect -860 -13452 -813 -9098
rect -749 -13452 -733 -9098
rect -461 -9209 -357 -8831
rect -141 -8942 -94 -4588
rect -30 -8942 -14 -4588
rect 258 -4699 362 -4321
rect 578 -4432 625 -78
rect 689 -4432 705 -78
rect 977 -189 1081 189
rect 1297 78 1344 4432
rect 1408 78 1424 4432
rect 1696 4321 1800 4699
rect 2016 4588 2063 8942
rect 2127 4588 2143 8942
rect 2415 8831 2519 9209
rect 2735 9098 2782 13452
rect 2846 9098 2862 13452
rect 2735 9082 2862 9098
rect 2735 8958 2839 9082
rect 2735 8942 2862 8958
rect 2306 8830 2628 8831
rect 2306 4700 2307 8830
rect 2627 4700 2628 8830
rect 2306 4699 2628 4700
rect 2016 4572 2143 4588
rect 2016 4448 2120 4572
rect 2016 4432 2143 4448
rect 1587 4320 1909 4321
rect 1587 190 1588 4320
rect 1908 190 1909 4320
rect 1587 189 1909 190
rect 1297 62 1424 78
rect 1297 -62 1401 62
rect 1297 -78 1424 -62
rect 868 -190 1190 -189
rect 868 -4320 869 -190
rect 1189 -4320 1190 -190
rect 868 -4321 1190 -4320
rect 578 -4448 705 -4432
rect 578 -4572 682 -4448
rect 578 -4588 705 -4572
rect 149 -4700 471 -4699
rect 149 -8830 150 -4700
rect 470 -8830 471 -4700
rect 149 -8831 471 -8830
rect -141 -8958 -14 -8942
rect -141 -9082 -37 -8958
rect -141 -9098 -14 -9082
rect -570 -9210 -248 -9209
rect -570 -13340 -569 -9210
rect -249 -13340 -248 -9210
rect -570 -13341 -248 -13340
rect -860 -13468 -733 -13452
rect -860 -13592 -756 -13468
rect -860 -13608 -733 -13592
rect -1289 -13720 -967 -13719
rect -1289 -17850 -1288 -13720
rect -968 -17850 -967 -13720
rect -1289 -17851 -967 -17850
rect -1579 -17978 -1452 -17962
rect -1579 -18102 -1475 -17978
rect -1579 -18118 -1452 -18102
rect -2008 -18230 -1686 -18229
rect -2008 -22360 -2007 -18230
rect -1687 -22360 -1686 -18230
rect -2008 -22361 -1686 -22360
rect -2298 -22488 -2171 -22472
rect -2298 -22612 -2194 -22488
rect -2298 -22628 -2171 -22612
rect -2727 -22740 -2405 -22739
rect -2727 -26870 -2726 -22740
rect -2406 -26870 -2405 -22740
rect -2727 -26871 -2405 -26870
rect -2618 -27249 -2514 -26871
rect -2298 -26982 -2251 -22628
rect -2187 -26982 -2171 -22628
rect -1899 -22739 -1795 -22361
rect -1579 -22472 -1532 -18118
rect -1468 -22472 -1452 -18118
rect -1180 -18229 -1076 -17851
rect -860 -17962 -813 -13608
rect -749 -17962 -733 -13608
rect -461 -13719 -357 -13341
rect -141 -13452 -94 -9098
rect -30 -13452 -14 -9098
rect 258 -9209 362 -8831
rect 578 -8942 625 -4588
rect 689 -8942 705 -4588
rect 977 -4699 1081 -4321
rect 1297 -4432 1344 -78
rect 1408 -4432 1424 -78
rect 1696 -189 1800 189
rect 2016 78 2063 4432
rect 2127 78 2143 4432
rect 2415 4321 2519 4699
rect 2735 4588 2782 8942
rect 2846 4588 2862 8942
rect 2735 4572 2862 4588
rect 2735 4448 2839 4572
rect 2735 4432 2862 4448
rect 2306 4320 2628 4321
rect 2306 190 2307 4320
rect 2627 190 2628 4320
rect 2306 189 2628 190
rect 2016 62 2143 78
rect 2016 -62 2120 62
rect 2016 -78 2143 -62
rect 1587 -190 1909 -189
rect 1587 -4320 1588 -190
rect 1908 -4320 1909 -190
rect 1587 -4321 1909 -4320
rect 1297 -4448 1424 -4432
rect 1297 -4572 1401 -4448
rect 1297 -4588 1424 -4572
rect 868 -4700 1190 -4699
rect 868 -8830 869 -4700
rect 1189 -8830 1190 -4700
rect 868 -8831 1190 -8830
rect 578 -8958 705 -8942
rect 578 -9082 682 -8958
rect 578 -9098 705 -9082
rect 149 -9210 471 -9209
rect 149 -13340 150 -9210
rect 470 -13340 471 -9210
rect 149 -13341 471 -13340
rect -141 -13468 -14 -13452
rect -141 -13592 -37 -13468
rect -141 -13608 -14 -13592
rect -570 -13720 -248 -13719
rect -570 -17850 -569 -13720
rect -249 -17850 -248 -13720
rect -570 -17851 -248 -17850
rect -860 -17978 -733 -17962
rect -860 -18102 -756 -17978
rect -860 -18118 -733 -18102
rect -1289 -18230 -967 -18229
rect -1289 -22360 -1288 -18230
rect -968 -22360 -967 -18230
rect -1289 -22361 -967 -22360
rect -1579 -22488 -1452 -22472
rect -1579 -22612 -1475 -22488
rect -1579 -22628 -1452 -22612
rect -2008 -22740 -1686 -22739
rect -2008 -26870 -2007 -22740
rect -1687 -26870 -1686 -22740
rect -2008 -26871 -1686 -26870
rect -2298 -26998 -2171 -26982
rect -2298 -27122 -2194 -26998
rect -2298 -27138 -2171 -27122
rect -2727 -27250 -2405 -27249
rect -2727 -31380 -2726 -27250
rect -2406 -31380 -2405 -27250
rect -2727 -31381 -2405 -31380
rect -2618 -31759 -2514 -31381
rect -2298 -31492 -2251 -27138
rect -2187 -31492 -2171 -27138
rect -1899 -27249 -1795 -26871
rect -1579 -26982 -1532 -22628
rect -1468 -26982 -1452 -22628
rect -1180 -22739 -1076 -22361
rect -860 -22472 -813 -18118
rect -749 -22472 -733 -18118
rect -461 -18229 -357 -17851
rect -141 -17962 -94 -13608
rect -30 -17962 -14 -13608
rect 258 -13719 362 -13341
rect 578 -13452 625 -9098
rect 689 -13452 705 -9098
rect 977 -9209 1081 -8831
rect 1297 -8942 1344 -4588
rect 1408 -8942 1424 -4588
rect 1696 -4699 1800 -4321
rect 2016 -4432 2063 -78
rect 2127 -4432 2143 -78
rect 2415 -189 2519 189
rect 2735 78 2782 4432
rect 2846 78 2862 4432
rect 2735 62 2862 78
rect 2735 -62 2839 62
rect 2735 -78 2862 -62
rect 2306 -190 2628 -189
rect 2306 -4320 2307 -190
rect 2627 -4320 2628 -190
rect 2306 -4321 2628 -4320
rect 2016 -4448 2143 -4432
rect 2016 -4572 2120 -4448
rect 2016 -4588 2143 -4572
rect 1587 -4700 1909 -4699
rect 1587 -8830 1588 -4700
rect 1908 -8830 1909 -4700
rect 1587 -8831 1909 -8830
rect 1297 -8958 1424 -8942
rect 1297 -9082 1401 -8958
rect 1297 -9098 1424 -9082
rect 868 -9210 1190 -9209
rect 868 -13340 869 -9210
rect 1189 -13340 1190 -9210
rect 868 -13341 1190 -13340
rect 578 -13468 705 -13452
rect 578 -13592 682 -13468
rect 578 -13608 705 -13592
rect 149 -13720 471 -13719
rect 149 -17850 150 -13720
rect 470 -17850 471 -13720
rect 149 -17851 471 -17850
rect -141 -17978 -14 -17962
rect -141 -18102 -37 -17978
rect -141 -18118 -14 -18102
rect -570 -18230 -248 -18229
rect -570 -22360 -569 -18230
rect -249 -22360 -248 -18230
rect -570 -22361 -248 -22360
rect -860 -22488 -733 -22472
rect -860 -22612 -756 -22488
rect -860 -22628 -733 -22612
rect -1289 -22740 -967 -22739
rect -1289 -26870 -1288 -22740
rect -968 -26870 -967 -22740
rect -1289 -26871 -967 -26870
rect -1579 -26998 -1452 -26982
rect -1579 -27122 -1475 -26998
rect -1579 -27138 -1452 -27122
rect -2008 -27250 -1686 -27249
rect -2008 -31380 -2007 -27250
rect -1687 -31380 -1686 -27250
rect -2008 -31381 -1686 -31380
rect -2298 -31508 -2171 -31492
rect -2298 -31632 -2194 -31508
rect -2298 -31648 -2171 -31632
rect -2727 -31760 -2405 -31759
rect -2727 -35890 -2726 -31760
rect -2406 -35890 -2405 -31760
rect -2727 -35891 -2405 -35890
rect -2618 -36080 -2514 -35891
rect -2298 -36002 -2251 -31648
rect -2187 -36002 -2171 -31648
rect -1899 -31759 -1795 -31381
rect -1579 -31492 -1532 -27138
rect -1468 -31492 -1452 -27138
rect -1180 -27249 -1076 -26871
rect -860 -26982 -813 -22628
rect -749 -26982 -733 -22628
rect -461 -22739 -357 -22361
rect -141 -22472 -94 -18118
rect -30 -22472 -14 -18118
rect 258 -18229 362 -17851
rect 578 -17962 625 -13608
rect 689 -17962 705 -13608
rect 977 -13719 1081 -13341
rect 1297 -13452 1344 -9098
rect 1408 -13452 1424 -9098
rect 1696 -9209 1800 -8831
rect 2016 -8942 2063 -4588
rect 2127 -8942 2143 -4588
rect 2415 -4699 2519 -4321
rect 2735 -4432 2782 -78
rect 2846 -4432 2862 -78
rect 2735 -4448 2862 -4432
rect 2735 -4572 2839 -4448
rect 2735 -4588 2862 -4572
rect 2306 -4700 2628 -4699
rect 2306 -8830 2307 -4700
rect 2627 -8830 2628 -4700
rect 2306 -8831 2628 -8830
rect 2016 -8958 2143 -8942
rect 2016 -9082 2120 -8958
rect 2016 -9098 2143 -9082
rect 1587 -9210 1909 -9209
rect 1587 -13340 1588 -9210
rect 1908 -13340 1909 -9210
rect 1587 -13341 1909 -13340
rect 1297 -13468 1424 -13452
rect 1297 -13592 1401 -13468
rect 1297 -13608 1424 -13592
rect 868 -13720 1190 -13719
rect 868 -17850 869 -13720
rect 1189 -17850 1190 -13720
rect 868 -17851 1190 -17850
rect 578 -17978 705 -17962
rect 578 -18102 682 -17978
rect 578 -18118 705 -18102
rect 149 -18230 471 -18229
rect 149 -22360 150 -18230
rect 470 -22360 471 -18230
rect 149 -22361 471 -22360
rect -141 -22488 -14 -22472
rect -141 -22612 -37 -22488
rect -141 -22628 -14 -22612
rect -570 -22740 -248 -22739
rect -570 -26870 -569 -22740
rect -249 -26870 -248 -22740
rect -570 -26871 -248 -26870
rect -860 -26998 -733 -26982
rect -860 -27122 -756 -26998
rect -860 -27138 -733 -27122
rect -1289 -27250 -967 -27249
rect -1289 -31380 -1288 -27250
rect -968 -31380 -967 -27250
rect -1289 -31381 -967 -31380
rect -1579 -31508 -1452 -31492
rect -1579 -31632 -1475 -31508
rect -1579 -31648 -1452 -31632
rect -2008 -31760 -1686 -31759
rect -2008 -35890 -2007 -31760
rect -1687 -35890 -1686 -31760
rect -2008 -35891 -1686 -35890
rect -2298 -36018 -2171 -36002
rect -2298 -36080 -2194 -36018
rect -1899 -36080 -1795 -35891
rect -1579 -36002 -1532 -31648
rect -1468 -36002 -1452 -31648
rect -1180 -31759 -1076 -31381
rect -860 -31492 -813 -27138
rect -749 -31492 -733 -27138
rect -461 -27249 -357 -26871
rect -141 -26982 -94 -22628
rect -30 -26982 -14 -22628
rect 258 -22739 362 -22361
rect 578 -22472 625 -18118
rect 689 -22472 705 -18118
rect 977 -18229 1081 -17851
rect 1297 -17962 1344 -13608
rect 1408 -17962 1424 -13608
rect 1696 -13719 1800 -13341
rect 2016 -13452 2063 -9098
rect 2127 -13452 2143 -9098
rect 2415 -9209 2519 -8831
rect 2735 -8942 2782 -4588
rect 2846 -8942 2862 -4588
rect 2735 -8958 2862 -8942
rect 2735 -9082 2839 -8958
rect 2735 -9098 2862 -9082
rect 2306 -9210 2628 -9209
rect 2306 -13340 2307 -9210
rect 2627 -13340 2628 -9210
rect 2306 -13341 2628 -13340
rect 2016 -13468 2143 -13452
rect 2016 -13592 2120 -13468
rect 2016 -13608 2143 -13592
rect 1587 -13720 1909 -13719
rect 1587 -17850 1588 -13720
rect 1908 -17850 1909 -13720
rect 1587 -17851 1909 -17850
rect 1297 -17978 1424 -17962
rect 1297 -18102 1401 -17978
rect 1297 -18118 1424 -18102
rect 868 -18230 1190 -18229
rect 868 -22360 869 -18230
rect 1189 -22360 1190 -18230
rect 868 -22361 1190 -22360
rect 578 -22488 705 -22472
rect 578 -22612 682 -22488
rect 578 -22628 705 -22612
rect 149 -22740 471 -22739
rect 149 -26870 150 -22740
rect 470 -26870 471 -22740
rect 149 -26871 471 -26870
rect -141 -26998 -14 -26982
rect -141 -27122 -37 -26998
rect -141 -27138 -14 -27122
rect -570 -27250 -248 -27249
rect -570 -31380 -569 -27250
rect -249 -31380 -248 -27250
rect -570 -31381 -248 -31380
rect -860 -31508 -733 -31492
rect -860 -31632 -756 -31508
rect -860 -31648 -733 -31632
rect -1289 -31760 -967 -31759
rect -1289 -35890 -1288 -31760
rect -968 -35890 -967 -31760
rect -1289 -35891 -967 -35890
rect -1579 -36018 -1452 -36002
rect -1579 -36080 -1475 -36018
rect -1180 -36080 -1076 -35891
rect -860 -36002 -813 -31648
rect -749 -36002 -733 -31648
rect -461 -31759 -357 -31381
rect -141 -31492 -94 -27138
rect -30 -31492 -14 -27138
rect 258 -27249 362 -26871
rect 578 -26982 625 -22628
rect 689 -26982 705 -22628
rect 977 -22739 1081 -22361
rect 1297 -22472 1344 -18118
rect 1408 -22472 1424 -18118
rect 1696 -18229 1800 -17851
rect 2016 -17962 2063 -13608
rect 2127 -17962 2143 -13608
rect 2415 -13719 2519 -13341
rect 2735 -13452 2782 -9098
rect 2846 -13452 2862 -9098
rect 2735 -13468 2862 -13452
rect 2735 -13592 2839 -13468
rect 2735 -13608 2862 -13592
rect 2306 -13720 2628 -13719
rect 2306 -17850 2307 -13720
rect 2627 -17850 2628 -13720
rect 2306 -17851 2628 -17850
rect 2016 -17978 2143 -17962
rect 2016 -18102 2120 -17978
rect 2016 -18118 2143 -18102
rect 1587 -18230 1909 -18229
rect 1587 -22360 1588 -18230
rect 1908 -22360 1909 -18230
rect 1587 -22361 1909 -22360
rect 1297 -22488 1424 -22472
rect 1297 -22612 1401 -22488
rect 1297 -22628 1424 -22612
rect 868 -22740 1190 -22739
rect 868 -26870 869 -22740
rect 1189 -26870 1190 -22740
rect 868 -26871 1190 -26870
rect 578 -26998 705 -26982
rect 578 -27122 682 -26998
rect 578 -27138 705 -27122
rect 149 -27250 471 -27249
rect 149 -31380 150 -27250
rect 470 -31380 471 -27250
rect 149 -31381 471 -31380
rect -141 -31508 -14 -31492
rect -141 -31632 -37 -31508
rect -141 -31648 -14 -31632
rect -570 -31760 -248 -31759
rect -570 -35890 -569 -31760
rect -249 -35890 -248 -31760
rect -570 -35891 -248 -35890
rect -860 -36018 -733 -36002
rect -860 -36080 -756 -36018
rect -461 -36080 -357 -35891
rect -141 -36002 -94 -31648
rect -30 -36002 -14 -31648
rect 258 -31759 362 -31381
rect 578 -31492 625 -27138
rect 689 -31492 705 -27138
rect 977 -27249 1081 -26871
rect 1297 -26982 1344 -22628
rect 1408 -26982 1424 -22628
rect 1696 -22739 1800 -22361
rect 2016 -22472 2063 -18118
rect 2127 -22472 2143 -18118
rect 2415 -18229 2519 -17851
rect 2735 -17962 2782 -13608
rect 2846 -17962 2862 -13608
rect 2735 -17978 2862 -17962
rect 2735 -18102 2839 -17978
rect 2735 -18118 2862 -18102
rect 2306 -18230 2628 -18229
rect 2306 -22360 2307 -18230
rect 2627 -22360 2628 -18230
rect 2306 -22361 2628 -22360
rect 2016 -22488 2143 -22472
rect 2016 -22612 2120 -22488
rect 2016 -22628 2143 -22612
rect 1587 -22740 1909 -22739
rect 1587 -26870 1588 -22740
rect 1908 -26870 1909 -22740
rect 1587 -26871 1909 -26870
rect 1297 -26998 1424 -26982
rect 1297 -27122 1401 -26998
rect 1297 -27138 1424 -27122
rect 868 -27250 1190 -27249
rect 868 -31380 869 -27250
rect 1189 -31380 1190 -27250
rect 868 -31381 1190 -31380
rect 578 -31508 705 -31492
rect 578 -31632 682 -31508
rect 578 -31648 705 -31632
rect 149 -31760 471 -31759
rect 149 -35890 150 -31760
rect 470 -35890 471 -31760
rect 149 -35891 471 -35890
rect -141 -36018 -14 -36002
rect -141 -36080 -37 -36018
rect 258 -36080 362 -35891
rect 578 -36002 625 -31648
rect 689 -36002 705 -31648
rect 977 -31759 1081 -31381
rect 1297 -31492 1344 -27138
rect 1408 -31492 1424 -27138
rect 1696 -27249 1800 -26871
rect 2016 -26982 2063 -22628
rect 2127 -26982 2143 -22628
rect 2415 -22739 2519 -22361
rect 2735 -22472 2782 -18118
rect 2846 -22472 2862 -18118
rect 2735 -22488 2862 -22472
rect 2735 -22612 2839 -22488
rect 2735 -22628 2862 -22612
rect 2306 -22740 2628 -22739
rect 2306 -26870 2307 -22740
rect 2627 -26870 2628 -22740
rect 2306 -26871 2628 -26870
rect 2016 -26998 2143 -26982
rect 2016 -27122 2120 -26998
rect 2016 -27138 2143 -27122
rect 1587 -27250 1909 -27249
rect 1587 -31380 1588 -27250
rect 1908 -31380 1909 -27250
rect 1587 -31381 1909 -31380
rect 1297 -31508 1424 -31492
rect 1297 -31632 1401 -31508
rect 1297 -31648 1424 -31632
rect 868 -31760 1190 -31759
rect 868 -35890 869 -31760
rect 1189 -35890 1190 -31760
rect 868 -35891 1190 -35890
rect 578 -36018 705 -36002
rect 578 -36080 682 -36018
rect 977 -36080 1081 -35891
rect 1297 -36002 1344 -31648
rect 1408 -36002 1424 -31648
rect 1696 -31759 1800 -31381
rect 2016 -31492 2063 -27138
rect 2127 -31492 2143 -27138
rect 2415 -27249 2519 -26871
rect 2735 -26982 2782 -22628
rect 2846 -26982 2862 -22628
rect 2735 -26998 2862 -26982
rect 2735 -27122 2839 -26998
rect 2735 -27138 2862 -27122
rect 2306 -27250 2628 -27249
rect 2306 -31380 2307 -27250
rect 2627 -31380 2628 -27250
rect 2306 -31381 2628 -31380
rect 2016 -31508 2143 -31492
rect 2016 -31632 2120 -31508
rect 2016 -31648 2143 -31632
rect 1587 -31760 1909 -31759
rect 1587 -35890 1588 -31760
rect 1908 -35890 1909 -31760
rect 1587 -35891 1909 -35890
rect 1297 -36018 1424 -36002
rect 1297 -36080 1401 -36018
rect 1696 -36080 1800 -35891
rect 2016 -36002 2063 -31648
rect 2127 -36002 2143 -31648
rect 2415 -31759 2519 -31381
rect 2735 -31492 2782 -27138
rect 2846 -31492 2862 -27138
rect 2735 -31508 2862 -31492
rect 2735 -31632 2839 -31508
rect 2735 -31648 2862 -31632
rect 2306 -31760 2628 -31759
rect 2306 -35890 2307 -31760
rect 2627 -35890 2628 -31760
rect 2306 -35891 2628 -35890
rect 2016 -36018 2143 -36002
rect 2016 -36080 2120 -36018
rect 2415 -36080 2519 -35891
rect 2735 -36002 2782 -31648
rect 2846 -36002 2862 -31648
rect 2735 -36018 2862 -36002
rect 2735 -36080 2839 -36018
<< properties >>
string FIXED_BBOX 2167 31620 2767 36030
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 8 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
