magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -386 72332 386 72360
rect -386 68098 302 72332
rect 366 68098 386 72332
rect -386 68070 386 68098
rect -386 67802 386 67830
rect -386 63568 302 67802
rect 366 63568 386 67802
rect -386 63540 386 63568
rect -386 63272 386 63300
rect -386 59038 302 63272
rect 366 59038 386 63272
rect -386 59010 386 59038
rect -386 58742 386 58770
rect -386 54508 302 58742
rect 366 54508 386 58742
rect -386 54480 386 54508
rect -386 54212 386 54240
rect -386 49978 302 54212
rect 366 49978 386 54212
rect -386 49950 386 49978
rect -386 49682 386 49710
rect -386 45448 302 49682
rect 366 45448 386 49682
rect -386 45420 386 45448
rect -386 45152 386 45180
rect -386 40918 302 45152
rect 366 40918 386 45152
rect -386 40890 386 40918
rect -386 40622 386 40650
rect -386 36388 302 40622
rect 366 36388 386 40622
rect -386 36360 386 36388
rect -386 36092 386 36120
rect -386 31858 302 36092
rect 366 31858 386 36092
rect -386 31830 386 31858
rect -386 31562 386 31590
rect -386 27328 302 31562
rect 366 27328 386 31562
rect -386 27300 386 27328
rect -386 27032 386 27060
rect -386 22798 302 27032
rect 366 22798 386 27032
rect -386 22770 386 22798
rect -386 22502 386 22530
rect -386 18268 302 22502
rect 366 18268 386 22502
rect -386 18240 386 18268
rect -386 17972 386 18000
rect -386 13738 302 17972
rect 366 13738 386 17972
rect -386 13710 386 13738
rect -386 13442 386 13470
rect -386 9208 302 13442
rect 366 9208 386 13442
rect -386 9180 386 9208
rect -386 8912 386 8940
rect -386 4678 302 8912
rect 366 4678 386 8912
rect -386 4650 386 4678
rect -386 4382 386 4410
rect -386 148 302 4382
rect 366 148 386 4382
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -4382 302 -148
rect 366 -4382 386 -148
rect -386 -4410 386 -4382
rect -386 -4678 386 -4650
rect -386 -8912 302 -4678
rect 366 -8912 386 -4678
rect -386 -8940 386 -8912
rect -386 -9208 386 -9180
rect -386 -13442 302 -9208
rect 366 -13442 386 -9208
rect -386 -13470 386 -13442
rect -386 -13738 386 -13710
rect -386 -17972 302 -13738
rect 366 -17972 386 -13738
rect -386 -18000 386 -17972
rect -386 -18268 386 -18240
rect -386 -22502 302 -18268
rect 366 -22502 386 -18268
rect -386 -22530 386 -22502
rect -386 -22798 386 -22770
rect -386 -27032 302 -22798
rect 366 -27032 386 -22798
rect -386 -27060 386 -27032
rect -386 -27328 386 -27300
rect -386 -31562 302 -27328
rect 366 -31562 386 -27328
rect -386 -31590 386 -31562
rect -386 -31858 386 -31830
rect -386 -36092 302 -31858
rect 366 -36092 386 -31858
rect -386 -36120 386 -36092
rect -386 -36388 386 -36360
rect -386 -40622 302 -36388
rect 366 -40622 386 -36388
rect -386 -40650 386 -40622
rect -386 -40918 386 -40890
rect -386 -45152 302 -40918
rect 366 -45152 386 -40918
rect -386 -45180 386 -45152
rect -386 -45448 386 -45420
rect -386 -49682 302 -45448
rect 366 -49682 386 -45448
rect -386 -49710 386 -49682
rect -386 -49978 386 -49950
rect -386 -54212 302 -49978
rect 366 -54212 386 -49978
rect -386 -54240 386 -54212
rect -386 -54508 386 -54480
rect -386 -58742 302 -54508
rect 366 -58742 386 -54508
rect -386 -58770 386 -58742
rect -386 -59038 386 -59010
rect -386 -63272 302 -59038
rect 366 -63272 386 -59038
rect -386 -63300 386 -63272
rect -386 -63568 386 -63540
rect -386 -67802 302 -63568
rect 366 -67802 386 -63568
rect -386 -67830 386 -67802
rect -386 -68098 386 -68070
rect -386 -72332 302 -68098
rect 366 -72332 386 -68098
rect -386 -72360 386 -72332
<< via3 >>
rect 302 68098 366 72332
rect 302 63568 366 67802
rect 302 59038 366 63272
rect 302 54508 366 58742
rect 302 49978 366 54212
rect 302 45448 366 49682
rect 302 40918 366 45152
rect 302 36388 366 40622
rect 302 31858 366 36092
rect 302 27328 366 31562
rect 302 22798 366 27032
rect 302 18268 366 22502
rect 302 13738 366 17972
rect 302 9208 366 13442
rect 302 4678 366 8912
rect 302 148 366 4382
rect 302 -4382 366 -148
rect 302 -8912 366 -4678
rect 302 -13442 366 -9208
rect 302 -17972 366 -13738
rect 302 -22502 366 -18268
rect 302 -27032 366 -22798
rect 302 -31562 366 -27328
rect 302 -36092 366 -31858
rect 302 -40622 366 -36388
rect 302 -45152 366 -40918
rect 302 -49682 366 -45448
rect 302 -54212 366 -49978
rect 302 -58742 366 -54508
rect 302 -63272 366 -59038
rect 302 -67802 366 -63568
rect 302 -72332 366 -68098
<< mimcap >>
rect -346 72280 54 72320
rect -346 68150 -306 72280
rect 14 68150 54 72280
rect -346 68110 54 68150
rect -346 67750 54 67790
rect -346 63620 -306 67750
rect 14 63620 54 67750
rect -346 63580 54 63620
rect -346 63220 54 63260
rect -346 59090 -306 63220
rect 14 59090 54 63220
rect -346 59050 54 59090
rect -346 58690 54 58730
rect -346 54560 -306 58690
rect 14 54560 54 58690
rect -346 54520 54 54560
rect -346 54160 54 54200
rect -346 50030 -306 54160
rect 14 50030 54 54160
rect -346 49990 54 50030
rect -346 49630 54 49670
rect -346 45500 -306 49630
rect 14 45500 54 49630
rect -346 45460 54 45500
rect -346 45100 54 45140
rect -346 40970 -306 45100
rect 14 40970 54 45100
rect -346 40930 54 40970
rect -346 40570 54 40610
rect -346 36440 -306 40570
rect 14 36440 54 40570
rect -346 36400 54 36440
rect -346 36040 54 36080
rect -346 31910 -306 36040
rect 14 31910 54 36040
rect -346 31870 54 31910
rect -346 31510 54 31550
rect -346 27380 -306 31510
rect 14 27380 54 31510
rect -346 27340 54 27380
rect -346 26980 54 27020
rect -346 22850 -306 26980
rect 14 22850 54 26980
rect -346 22810 54 22850
rect -346 22450 54 22490
rect -346 18320 -306 22450
rect 14 18320 54 22450
rect -346 18280 54 18320
rect -346 17920 54 17960
rect -346 13790 -306 17920
rect 14 13790 54 17920
rect -346 13750 54 13790
rect -346 13390 54 13430
rect -346 9260 -306 13390
rect 14 9260 54 13390
rect -346 9220 54 9260
rect -346 8860 54 8900
rect -346 4730 -306 8860
rect 14 4730 54 8860
rect -346 4690 54 4730
rect -346 4330 54 4370
rect -346 200 -306 4330
rect 14 200 54 4330
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -4330 -306 -200
rect 14 -4330 54 -200
rect -346 -4370 54 -4330
rect -346 -4730 54 -4690
rect -346 -8860 -306 -4730
rect 14 -8860 54 -4730
rect -346 -8900 54 -8860
rect -346 -9260 54 -9220
rect -346 -13390 -306 -9260
rect 14 -13390 54 -9260
rect -346 -13430 54 -13390
rect -346 -13790 54 -13750
rect -346 -17920 -306 -13790
rect 14 -17920 54 -13790
rect -346 -17960 54 -17920
rect -346 -18320 54 -18280
rect -346 -22450 -306 -18320
rect 14 -22450 54 -18320
rect -346 -22490 54 -22450
rect -346 -22850 54 -22810
rect -346 -26980 -306 -22850
rect 14 -26980 54 -22850
rect -346 -27020 54 -26980
rect -346 -27380 54 -27340
rect -346 -31510 -306 -27380
rect 14 -31510 54 -27380
rect -346 -31550 54 -31510
rect -346 -31910 54 -31870
rect -346 -36040 -306 -31910
rect 14 -36040 54 -31910
rect -346 -36080 54 -36040
rect -346 -36440 54 -36400
rect -346 -40570 -306 -36440
rect 14 -40570 54 -36440
rect -346 -40610 54 -40570
rect -346 -40970 54 -40930
rect -346 -45100 -306 -40970
rect 14 -45100 54 -40970
rect -346 -45140 54 -45100
rect -346 -45500 54 -45460
rect -346 -49630 -306 -45500
rect 14 -49630 54 -45500
rect -346 -49670 54 -49630
rect -346 -50030 54 -49990
rect -346 -54160 -306 -50030
rect 14 -54160 54 -50030
rect -346 -54200 54 -54160
rect -346 -54560 54 -54520
rect -346 -58690 -306 -54560
rect 14 -58690 54 -54560
rect -346 -58730 54 -58690
rect -346 -59090 54 -59050
rect -346 -63220 -306 -59090
rect 14 -63220 54 -59090
rect -346 -63260 54 -63220
rect -346 -63620 54 -63580
rect -346 -67750 -306 -63620
rect 14 -67750 54 -63620
rect -346 -67790 54 -67750
rect -346 -68150 54 -68110
rect -346 -72280 -306 -68150
rect 14 -72280 54 -68150
rect -346 -72320 54 -72280
<< mimcapcontact >>
rect -306 68150 14 72280
rect -306 63620 14 67750
rect -306 59090 14 63220
rect -306 54560 14 58690
rect -306 50030 14 54160
rect -306 45500 14 49630
rect -306 40970 14 45100
rect -306 36440 14 40570
rect -306 31910 14 36040
rect -306 27380 14 31510
rect -306 22850 14 26980
rect -306 18320 14 22450
rect -306 13790 14 17920
rect -306 9260 14 13390
rect -306 4730 14 8860
rect -306 200 14 4330
rect -306 -4330 14 -200
rect -306 -8860 14 -4730
rect -306 -13390 14 -9260
rect -306 -17920 14 -13790
rect -306 -22450 14 -18320
rect -306 -26980 14 -22850
rect -306 -31510 14 -27380
rect -306 -36040 14 -31910
rect -306 -40570 14 -36440
rect -306 -45100 14 -40970
rect -306 -49630 14 -45500
rect -306 -54160 14 -50030
rect -306 -58690 14 -54560
rect -306 -63220 14 -59090
rect -306 -67750 14 -63620
rect -306 -72280 14 -68150
<< metal4 >>
rect -198 72281 -94 72480
rect 282 72332 386 72480
rect -307 72280 15 72281
rect -307 68150 -306 72280
rect 14 68150 15 72280
rect -307 68149 15 68150
rect -198 67751 -94 68149
rect 282 68098 302 72332
rect 366 68098 386 72332
rect 282 67802 386 68098
rect -307 67750 15 67751
rect -307 63620 -306 67750
rect 14 63620 15 67750
rect -307 63619 15 63620
rect -198 63221 -94 63619
rect 282 63568 302 67802
rect 366 63568 386 67802
rect 282 63272 386 63568
rect -307 63220 15 63221
rect -307 59090 -306 63220
rect 14 59090 15 63220
rect -307 59089 15 59090
rect -198 58691 -94 59089
rect 282 59038 302 63272
rect 366 59038 386 63272
rect 282 58742 386 59038
rect -307 58690 15 58691
rect -307 54560 -306 58690
rect 14 54560 15 58690
rect -307 54559 15 54560
rect -198 54161 -94 54559
rect 282 54508 302 58742
rect 366 54508 386 58742
rect 282 54212 386 54508
rect -307 54160 15 54161
rect -307 50030 -306 54160
rect 14 50030 15 54160
rect -307 50029 15 50030
rect -198 49631 -94 50029
rect 282 49978 302 54212
rect 366 49978 386 54212
rect 282 49682 386 49978
rect -307 49630 15 49631
rect -307 45500 -306 49630
rect 14 45500 15 49630
rect -307 45499 15 45500
rect -198 45101 -94 45499
rect 282 45448 302 49682
rect 366 45448 386 49682
rect 282 45152 386 45448
rect -307 45100 15 45101
rect -307 40970 -306 45100
rect 14 40970 15 45100
rect -307 40969 15 40970
rect -198 40571 -94 40969
rect 282 40918 302 45152
rect 366 40918 386 45152
rect 282 40622 386 40918
rect -307 40570 15 40571
rect -307 36440 -306 40570
rect 14 36440 15 40570
rect -307 36439 15 36440
rect -198 36041 -94 36439
rect 282 36388 302 40622
rect 366 36388 386 40622
rect 282 36092 386 36388
rect -307 36040 15 36041
rect -307 31910 -306 36040
rect 14 31910 15 36040
rect -307 31909 15 31910
rect -198 31511 -94 31909
rect 282 31858 302 36092
rect 366 31858 386 36092
rect 282 31562 386 31858
rect -307 31510 15 31511
rect -307 27380 -306 31510
rect 14 27380 15 31510
rect -307 27379 15 27380
rect -198 26981 -94 27379
rect 282 27328 302 31562
rect 366 27328 386 31562
rect 282 27032 386 27328
rect -307 26980 15 26981
rect -307 22850 -306 26980
rect 14 22850 15 26980
rect -307 22849 15 22850
rect -198 22451 -94 22849
rect 282 22798 302 27032
rect 366 22798 386 27032
rect 282 22502 386 22798
rect -307 22450 15 22451
rect -307 18320 -306 22450
rect 14 18320 15 22450
rect -307 18319 15 18320
rect -198 17921 -94 18319
rect 282 18268 302 22502
rect 366 18268 386 22502
rect 282 17972 386 18268
rect -307 17920 15 17921
rect -307 13790 -306 17920
rect 14 13790 15 17920
rect -307 13789 15 13790
rect -198 13391 -94 13789
rect 282 13738 302 17972
rect 366 13738 386 17972
rect 282 13442 386 13738
rect -307 13390 15 13391
rect -307 9260 -306 13390
rect 14 9260 15 13390
rect -307 9259 15 9260
rect -198 8861 -94 9259
rect 282 9208 302 13442
rect 366 9208 386 13442
rect 282 8912 386 9208
rect -307 8860 15 8861
rect -307 4730 -306 8860
rect 14 4730 15 8860
rect -307 4729 15 4730
rect -198 4331 -94 4729
rect 282 4678 302 8912
rect 366 4678 386 8912
rect 282 4382 386 4678
rect -307 4330 15 4331
rect -307 200 -306 4330
rect 14 200 15 4330
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 4382
rect 366 148 386 4382
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -4330 -306 -200
rect 14 -4330 15 -200
rect -307 -4331 15 -4330
rect -198 -4729 -94 -4331
rect 282 -4382 302 -148
rect 366 -4382 386 -148
rect 282 -4678 386 -4382
rect -307 -4730 15 -4729
rect -307 -8860 -306 -4730
rect 14 -8860 15 -4730
rect -307 -8861 15 -8860
rect -198 -9259 -94 -8861
rect 282 -8912 302 -4678
rect 366 -8912 386 -4678
rect 282 -9208 386 -8912
rect -307 -9260 15 -9259
rect -307 -13390 -306 -9260
rect 14 -13390 15 -9260
rect -307 -13391 15 -13390
rect -198 -13789 -94 -13391
rect 282 -13442 302 -9208
rect 366 -13442 386 -9208
rect 282 -13738 386 -13442
rect -307 -13790 15 -13789
rect -307 -17920 -306 -13790
rect 14 -17920 15 -13790
rect -307 -17921 15 -17920
rect -198 -18319 -94 -17921
rect 282 -17972 302 -13738
rect 366 -17972 386 -13738
rect 282 -18268 386 -17972
rect -307 -18320 15 -18319
rect -307 -22450 -306 -18320
rect 14 -22450 15 -18320
rect -307 -22451 15 -22450
rect -198 -22849 -94 -22451
rect 282 -22502 302 -18268
rect 366 -22502 386 -18268
rect 282 -22798 386 -22502
rect -307 -22850 15 -22849
rect -307 -26980 -306 -22850
rect 14 -26980 15 -22850
rect -307 -26981 15 -26980
rect -198 -27379 -94 -26981
rect 282 -27032 302 -22798
rect 366 -27032 386 -22798
rect 282 -27328 386 -27032
rect -307 -27380 15 -27379
rect -307 -31510 -306 -27380
rect 14 -31510 15 -27380
rect -307 -31511 15 -31510
rect -198 -31909 -94 -31511
rect 282 -31562 302 -27328
rect 366 -31562 386 -27328
rect 282 -31858 386 -31562
rect -307 -31910 15 -31909
rect -307 -36040 -306 -31910
rect 14 -36040 15 -31910
rect -307 -36041 15 -36040
rect -198 -36439 -94 -36041
rect 282 -36092 302 -31858
rect 366 -36092 386 -31858
rect 282 -36388 386 -36092
rect -307 -36440 15 -36439
rect -307 -40570 -306 -36440
rect 14 -40570 15 -36440
rect -307 -40571 15 -40570
rect -198 -40969 -94 -40571
rect 282 -40622 302 -36388
rect 366 -40622 386 -36388
rect 282 -40918 386 -40622
rect -307 -40970 15 -40969
rect -307 -45100 -306 -40970
rect 14 -45100 15 -40970
rect -307 -45101 15 -45100
rect -198 -45499 -94 -45101
rect 282 -45152 302 -40918
rect 366 -45152 386 -40918
rect 282 -45448 386 -45152
rect -307 -45500 15 -45499
rect -307 -49630 -306 -45500
rect 14 -49630 15 -45500
rect -307 -49631 15 -49630
rect -198 -50029 -94 -49631
rect 282 -49682 302 -45448
rect 366 -49682 386 -45448
rect 282 -49978 386 -49682
rect -307 -50030 15 -50029
rect -307 -54160 -306 -50030
rect 14 -54160 15 -50030
rect -307 -54161 15 -54160
rect -198 -54559 -94 -54161
rect 282 -54212 302 -49978
rect 366 -54212 386 -49978
rect 282 -54508 386 -54212
rect -307 -54560 15 -54559
rect -307 -58690 -306 -54560
rect 14 -58690 15 -54560
rect -307 -58691 15 -58690
rect -198 -59089 -94 -58691
rect 282 -58742 302 -54508
rect 366 -58742 386 -54508
rect 282 -59038 386 -58742
rect -307 -59090 15 -59089
rect -307 -63220 -306 -59090
rect 14 -63220 15 -59090
rect -307 -63221 15 -63220
rect -198 -63619 -94 -63221
rect 282 -63272 302 -59038
rect 366 -63272 386 -59038
rect 282 -63568 386 -63272
rect -307 -63620 15 -63619
rect -307 -67750 -306 -63620
rect 14 -67750 15 -63620
rect -307 -67751 15 -67750
rect -198 -68149 -94 -67751
rect 282 -67802 302 -63568
rect 366 -67802 386 -63568
rect 282 -68098 386 -67802
rect -307 -68150 15 -68149
rect -307 -72280 -306 -68150
rect 14 -72280 15 -68150
rect -307 -72281 15 -72280
rect -198 -72480 -94 -72281
rect 282 -72332 302 -68098
rect 366 -72332 386 -68098
rect 282 -72480 386 -72332
<< properties >>
string FIXED_BBOX -386 68070 94 72360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 1 ny 32 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
