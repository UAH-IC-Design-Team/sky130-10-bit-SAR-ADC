magic
tech sky130A
magscale 1 2
timestamp 1666291486
<< metal4 >>
rect -2796 1039 -1698 1080
rect -2796 561 -1954 1039
rect -1718 561 -1698 1039
rect -2796 520 -1698 561
rect -1298 1039 -200 1080
rect -1298 561 -456 1039
rect -220 561 -200 1039
rect -1298 520 -200 561
rect 200 1039 1298 1080
rect 200 561 1042 1039
rect 1278 561 1298 1039
rect 200 520 1298 561
rect 1698 1039 2796 1080
rect 1698 561 2540 1039
rect 2776 561 2796 1039
rect 1698 520 2796 561
rect -2796 239 -1698 280
rect -2796 -239 -1954 239
rect -1718 -239 -1698 239
rect -2796 -280 -1698 -239
rect -1298 239 -200 280
rect -1298 -239 -456 239
rect -220 -239 -200 239
rect -1298 -280 -200 -239
rect 200 239 1298 280
rect 200 -239 1042 239
rect 1278 -239 1298 239
rect 200 -280 1298 -239
rect 1698 239 2796 280
rect 1698 -239 2540 239
rect 2776 -239 2796 239
rect 1698 -280 2796 -239
rect -2796 -561 -1698 -520
rect -2796 -1039 -1954 -561
rect -1718 -1039 -1698 -561
rect -2796 -1080 -1698 -1039
rect -1298 -561 -200 -520
rect -1298 -1039 -456 -561
rect -220 -1039 -200 -561
rect -1298 -1080 -200 -1039
rect 200 -561 1298 -520
rect 200 -1039 1042 -561
rect 1278 -1039 1298 -561
rect 200 -1080 1298 -1039
rect 1698 -561 2796 -520
rect 1698 -1039 2540 -561
rect 2776 -1039 2796 -561
rect 1698 -1080 2796 -1039
<< via4 >>
rect -1954 561 -1718 1039
rect -456 561 -220 1039
rect 1042 561 1278 1039
rect 2540 561 2776 1039
rect -1954 -239 -1718 239
rect -456 -239 -220 239
rect 1042 -239 1278 239
rect 2540 -239 2776 239
rect -1954 -1039 -1718 -561
rect -456 -1039 -220 -561
rect 1042 -1039 1278 -561
rect 2540 -1039 2776 -561
<< mimcap2 >>
rect -2716 960 -2316 1000
rect -2716 640 -2676 960
rect -2356 640 -2316 960
rect -2716 600 -2316 640
rect -1218 960 -818 1000
rect -1218 640 -1178 960
rect -858 640 -818 960
rect -1218 600 -818 640
rect 280 960 680 1000
rect 280 640 320 960
rect 640 640 680 960
rect 280 600 680 640
rect 1778 960 2178 1000
rect 1778 640 1818 960
rect 2138 640 2178 960
rect 1778 600 2178 640
rect -2716 160 -2316 200
rect -2716 -160 -2676 160
rect -2356 -160 -2316 160
rect -2716 -200 -2316 -160
rect -1218 160 -818 200
rect -1218 -160 -1178 160
rect -858 -160 -818 160
rect -1218 -200 -818 -160
rect 280 160 680 200
rect 280 -160 320 160
rect 640 -160 680 160
rect 280 -200 680 -160
rect 1778 160 2178 200
rect 1778 -160 1818 160
rect 2138 -160 2178 160
rect 1778 -200 2178 -160
rect -2716 -640 -2316 -600
rect -2716 -960 -2676 -640
rect -2356 -960 -2316 -640
rect -2716 -1000 -2316 -960
rect -1218 -640 -818 -600
rect -1218 -960 -1178 -640
rect -858 -960 -818 -640
rect -1218 -1000 -818 -960
rect 280 -640 680 -600
rect 280 -960 320 -640
rect 640 -960 680 -640
rect 280 -1000 680 -960
rect 1778 -640 2178 -600
rect 1778 -960 1818 -640
rect 2138 -960 2178 -640
rect 1778 -1000 2178 -960
<< mimcap2contact >>
rect -2676 640 -2356 960
rect -1178 640 -858 960
rect 320 640 640 960
rect 1818 640 2138 960
rect -2676 -160 -2356 160
rect -1178 -160 -858 160
rect 320 -160 640 160
rect 1818 -160 2138 160
rect -2676 -960 -2356 -640
rect -1178 -960 -858 -640
rect 320 -960 640 -640
rect 1818 -960 2138 -640
<< metal5 >>
rect -2676 984 -2356 1200
rect -1996 1039 -1676 1200
rect -2700 960 -2332 984
rect -2700 640 -2676 960
rect -2356 640 -2332 960
rect -2700 616 -2332 640
rect -2676 184 -2356 616
rect -1996 561 -1954 1039
rect -1718 561 -1676 1039
rect -1178 984 -858 1200
rect -498 1039 -178 1200
rect -1202 960 -834 984
rect -1202 640 -1178 960
rect -858 640 -834 960
rect -1202 616 -834 640
rect -1996 239 -1676 561
rect -2700 160 -2332 184
rect -2700 -160 -2676 160
rect -2356 -160 -2332 160
rect -2700 -184 -2332 -160
rect -2676 -616 -2356 -184
rect -1996 -239 -1954 239
rect -1718 -239 -1676 239
rect -1178 184 -858 616
rect -498 561 -456 1039
rect -220 561 -178 1039
rect 320 984 640 1200
rect 1000 1039 1320 1200
rect 296 960 664 984
rect 296 640 320 960
rect 640 640 664 960
rect 296 616 664 640
rect -498 239 -178 561
rect -1202 160 -834 184
rect -1202 -160 -1178 160
rect -858 -160 -834 160
rect -1202 -184 -834 -160
rect -1996 -561 -1676 -239
rect -2700 -640 -2332 -616
rect -2700 -960 -2676 -640
rect -2356 -960 -2332 -640
rect -2700 -984 -2332 -960
rect -2676 -1200 -2356 -984
rect -1996 -1039 -1954 -561
rect -1718 -1039 -1676 -561
rect -1178 -616 -858 -184
rect -498 -239 -456 239
rect -220 -239 -178 239
rect 320 184 640 616
rect 1000 561 1042 1039
rect 1278 561 1320 1039
rect 1818 984 2138 1200
rect 2498 1039 2818 1200
rect 1794 960 2162 984
rect 1794 640 1818 960
rect 2138 640 2162 960
rect 1794 616 2162 640
rect 1000 239 1320 561
rect 296 160 664 184
rect 296 -160 320 160
rect 640 -160 664 160
rect 296 -184 664 -160
rect -498 -561 -178 -239
rect -1202 -640 -834 -616
rect -1202 -960 -1178 -640
rect -858 -960 -834 -640
rect -1202 -984 -834 -960
rect -1996 -1200 -1676 -1039
rect -1178 -1200 -858 -984
rect -498 -1039 -456 -561
rect -220 -1039 -178 -561
rect 320 -616 640 -184
rect 1000 -239 1042 239
rect 1278 -239 1320 239
rect 1818 184 2138 616
rect 2498 561 2540 1039
rect 2776 561 2818 1039
rect 2498 239 2818 561
rect 1794 160 2162 184
rect 1794 -160 1818 160
rect 2138 -160 2162 160
rect 1794 -184 2162 -160
rect 1000 -561 1320 -239
rect 296 -640 664 -616
rect 296 -960 320 -640
rect 640 -960 664 -640
rect 296 -984 664 -960
rect -498 -1200 -178 -1039
rect 320 -1200 640 -984
rect 1000 -1039 1042 -561
rect 1278 -1039 1320 -561
rect 1818 -616 2138 -184
rect 2498 -239 2540 239
rect 2776 -239 2818 239
rect 2498 -561 2818 -239
rect 1794 -640 2162 -616
rect 1794 -960 1818 -640
rect 2138 -960 2162 -640
rect 1794 -984 2162 -960
rect 1000 -1200 1320 -1039
rect 1818 -1200 2138 -984
rect 2498 -1039 2540 -561
rect 2776 -1039 2818 -561
rect 2498 -1200 2818 -1039
<< properties >>
string FIXED_BBOX 1698 520 2258 1080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 4 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
