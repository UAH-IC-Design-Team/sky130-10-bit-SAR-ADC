magic
tech sky130A
magscale 1 2
timestamp 1666552007
<< error_p >>
rect -29 763 29 769
rect -29 729 -17 763
rect -29 723 29 729
rect -29 471 29 477
rect -29 437 -17 471
rect -29 431 29 437
rect -29 363 29 369
rect -29 329 -17 363
rect -29 323 29 329
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -329 29 -323
rect -29 -363 -17 -329
rect -29 -369 29 -363
rect -29 -437 29 -431
rect -29 -471 -17 -437
rect -29 -477 29 -471
rect -29 -729 29 -723
rect -29 -763 -17 -729
rect -29 -769 29 -763
<< pwell >>
rect -211 -901 211 901
<< nmos >>
rect -15 509 15 691
rect -15 109 15 291
rect -15 -291 15 -109
rect -15 -691 15 -509
<< ndiff >>
rect -73 679 -15 691
rect -73 521 -61 679
rect -27 521 -15 679
rect -73 509 -15 521
rect 15 679 73 691
rect 15 521 27 679
rect 61 521 73 679
rect 15 509 73 521
rect -73 279 -15 291
rect -73 121 -61 279
rect -27 121 -15 279
rect -73 109 -15 121
rect 15 279 73 291
rect 15 121 27 279
rect 61 121 73 279
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -279 -61 -121
rect -27 -279 -15 -121
rect -73 -291 -15 -279
rect 15 -121 73 -109
rect 15 -279 27 -121
rect 61 -279 73 -121
rect 15 -291 73 -279
rect -73 -521 -15 -509
rect -73 -679 -61 -521
rect -27 -679 -15 -521
rect -73 -691 -15 -679
rect 15 -521 73 -509
rect 15 -679 27 -521
rect 61 -679 73 -521
rect 15 -691 73 -679
<< ndiffc >>
rect -61 521 -27 679
rect 27 521 61 679
rect -61 121 -27 279
rect 27 121 61 279
rect -61 -279 -27 -121
rect 27 -279 61 -121
rect -61 -679 -27 -521
rect 27 -679 61 -521
<< psubdiff >>
rect -175 831 -79 865
rect 79 831 175 865
rect -175 -831 -141 831
rect 141 769 175 831
rect 141 -831 175 -769
rect -175 -865 -79 -831
rect 79 -865 175 -831
<< psubdiffcont >>
rect -79 831 79 865
rect 141 -769 175 769
rect -79 -865 79 -831
<< poly >>
rect -33 763 33 779
rect -33 729 -17 763
rect 17 729 33 763
rect -33 713 33 729
rect -15 691 15 713
rect -15 487 15 509
rect -33 471 33 487
rect -33 437 -17 471
rect 17 437 33 471
rect -33 421 33 437
rect -33 363 33 379
rect -33 329 -17 363
rect 17 329 33 363
rect -33 313 33 329
rect -15 291 15 313
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -313 15 -291
rect -33 -329 33 -313
rect -33 -363 -17 -329
rect 17 -363 33 -329
rect -33 -379 33 -363
rect -33 -437 33 -421
rect -33 -471 -17 -437
rect 17 -471 33 -437
rect -33 -487 33 -471
rect -15 -509 15 -487
rect -15 -713 15 -691
rect -33 -729 33 -713
rect -33 -763 -17 -729
rect 17 -763 33 -729
rect -33 -779 33 -763
<< polycont >>
rect -17 729 17 763
rect -17 437 17 471
rect -17 329 17 363
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -363 17 -329
rect -17 -471 17 -437
rect -17 -763 17 -729
<< locali >>
rect -95 831 -79 865
rect 79 831 95 865
rect 141 769 175 785
rect -33 729 -17 763
rect 17 729 33 763
rect -61 679 -27 695
rect -61 505 -27 521
rect 27 679 61 695
rect 27 505 61 521
rect -33 437 -17 471
rect 17 437 33 471
rect -33 329 -17 363
rect 17 329 33 363
rect -61 279 -27 295
rect -61 105 -27 121
rect 27 279 61 295
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -295 -27 -279
rect 27 -121 61 -105
rect 27 -295 61 -279
rect -33 -363 -17 -329
rect 17 -363 33 -329
rect -33 -471 -17 -437
rect 17 -471 33 -437
rect -61 -521 -27 -505
rect -61 -695 -27 -679
rect 27 -521 61 -505
rect 27 -695 61 -679
rect -33 -763 -17 -729
rect 17 -763 33 -729
rect 141 -785 175 -769
rect -95 -865 -79 -831
rect 79 -865 95 -831
<< viali >>
rect -17 729 17 763
rect -61 521 -27 679
rect 27 521 61 679
rect -17 437 17 471
rect -17 329 17 363
rect -61 121 -27 279
rect 27 121 61 279
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -279 -27 -121
rect 27 -279 61 -121
rect -17 -363 17 -329
rect -17 -471 17 -437
rect -61 -679 -27 -521
rect 27 -679 61 -521
rect -17 -763 17 -729
<< metal1 >>
rect -29 763 29 769
rect -29 729 -17 763
rect 17 729 29 763
rect -29 723 29 729
rect -67 679 -21 691
rect -67 521 -61 679
rect -27 521 -21 679
rect -67 509 -21 521
rect 21 679 67 691
rect 21 521 27 679
rect 61 521 67 679
rect 21 509 67 521
rect -29 471 29 477
rect -29 437 -17 471
rect 17 437 29 471
rect -29 431 29 437
rect -29 363 29 369
rect -29 329 -17 363
rect 17 329 29 363
rect -29 323 29 329
rect -67 279 -21 291
rect -67 121 -61 279
rect -27 121 -21 279
rect -67 109 -21 121
rect 21 279 67 291
rect 21 121 27 279
rect 61 121 67 279
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -279 -61 -121
rect -27 -279 -21 -121
rect -67 -291 -21 -279
rect 21 -121 67 -109
rect 21 -279 27 -121
rect 61 -279 67 -121
rect 21 -291 67 -279
rect -29 -329 29 -323
rect -29 -363 -17 -329
rect 17 -363 29 -329
rect -29 -369 29 -363
rect -29 -437 29 -431
rect -29 -471 -17 -437
rect 17 -471 29 -437
rect -29 -477 29 -471
rect -67 -521 -21 -509
rect -67 -679 -61 -521
rect -27 -679 -21 -521
rect -67 -691 -21 -679
rect 21 -521 67 -509
rect 21 -679 27 -521
rect 61 -679 67 -521
rect 21 -691 67 -679
rect -29 -729 29 -723
rect -29 -763 -17 -729
rect 17 -763 29 -729
rect -29 -769 29 -763
<< properties >>
string FIXED_BBOX -158 -848 158 848
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
