magic
tech sky130A
magscale 1 2
timestamp 1666918349
<< error_p >>
rect -29 6053 29 6059
rect -29 6019 -17 6053
rect -29 6013 29 6019
rect -29 4943 29 4949
rect -29 4909 -17 4943
rect -29 4903 29 4909
rect -29 4835 29 4841
rect -29 4801 -17 4835
rect -29 4795 29 4801
rect -29 3725 29 3731
rect -29 3691 -17 3725
rect -29 3685 29 3691
rect -29 3617 29 3623
rect -29 3583 -17 3617
rect -29 3577 29 3583
rect -29 2507 29 2513
rect -29 2473 -17 2507
rect -29 2467 29 2473
rect -29 2399 29 2405
rect -29 2365 -17 2399
rect -29 2359 29 2365
rect -29 1289 29 1295
rect -29 1255 -17 1289
rect -29 1249 29 1255
rect -29 1181 29 1187
rect -29 1147 -17 1181
rect -29 1141 29 1147
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -1147 29 -1141
rect -29 -1181 -17 -1147
rect -29 -1187 29 -1181
rect -29 -1255 29 -1249
rect -29 -1289 -17 -1255
rect -29 -1295 29 -1289
rect -29 -2365 29 -2359
rect -29 -2399 -17 -2365
rect -29 -2405 29 -2399
rect -29 -2473 29 -2467
rect -29 -2507 -17 -2473
rect -29 -2513 29 -2507
rect -29 -3583 29 -3577
rect -29 -3617 -17 -3583
rect -29 -3623 29 -3617
rect -29 -3691 29 -3685
rect -29 -3725 -17 -3691
rect -29 -3731 29 -3725
rect -29 -4801 29 -4795
rect -29 -4835 -17 -4801
rect -29 -4841 29 -4835
rect -29 -4909 29 -4903
rect -29 -4943 -17 -4909
rect -29 -4949 29 -4943
rect -29 -6019 29 -6013
rect -29 -6053 -17 -6019
rect -29 -6059 29 -6053
<< pwell >>
rect -211 -6191 211 6191
<< nmos >>
rect -15 4981 15 5981
rect -15 3763 15 4763
rect -15 2545 15 3545
rect -15 1327 15 2327
rect -15 109 15 1109
rect -15 -1109 15 -109
rect -15 -2327 15 -1327
rect -15 -3545 15 -2545
rect -15 -4763 15 -3763
rect -15 -5981 15 -4981
<< ndiff >>
rect -73 5969 -15 5981
rect -73 4993 -61 5969
rect -27 4993 -15 5969
rect -73 4981 -15 4993
rect 15 5969 73 5981
rect 15 4993 27 5969
rect 61 4993 73 5969
rect 15 4981 73 4993
rect -73 4751 -15 4763
rect -73 3775 -61 4751
rect -27 3775 -15 4751
rect -73 3763 -15 3775
rect 15 4751 73 4763
rect 15 3775 27 4751
rect 61 3775 73 4751
rect 15 3763 73 3775
rect -73 3533 -15 3545
rect -73 2557 -61 3533
rect -27 2557 -15 3533
rect -73 2545 -15 2557
rect 15 3533 73 3545
rect 15 2557 27 3533
rect 61 2557 73 3533
rect 15 2545 73 2557
rect -73 2315 -15 2327
rect -73 1339 -61 2315
rect -27 1339 -15 2315
rect -73 1327 -15 1339
rect 15 2315 73 2327
rect 15 1339 27 2315
rect 61 1339 73 2315
rect 15 1327 73 1339
rect -73 1097 -15 1109
rect -73 121 -61 1097
rect -27 121 -15 1097
rect -73 109 -15 121
rect 15 1097 73 1109
rect 15 121 27 1097
rect 61 121 73 1097
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -1097 -61 -121
rect -27 -1097 -15 -121
rect -73 -1109 -15 -1097
rect 15 -121 73 -109
rect 15 -1097 27 -121
rect 61 -1097 73 -121
rect 15 -1109 73 -1097
rect -73 -1339 -15 -1327
rect -73 -2315 -61 -1339
rect -27 -2315 -15 -1339
rect -73 -2327 -15 -2315
rect 15 -1339 73 -1327
rect 15 -2315 27 -1339
rect 61 -2315 73 -1339
rect 15 -2327 73 -2315
rect -73 -2557 -15 -2545
rect -73 -3533 -61 -2557
rect -27 -3533 -15 -2557
rect -73 -3545 -15 -3533
rect 15 -2557 73 -2545
rect 15 -3533 27 -2557
rect 61 -3533 73 -2557
rect 15 -3545 73 -3533
rect -73 -3775 -15 -3763
rect -73 -4751 -61 -3775
rect -27 -4751 -15 -3775
rect -73 -4763 -15 -4751
rect 15 -3775 73 -3763
rect 15 -4751 27 -3775
rect 61 -4751 73 -3775
rect 15 -4763 73 -4751
rect -73 -4993 -15 -4981
rect -73 -5969 -61 -4993
rect -27 -5969 -15 -4993
rect -73 -5981 -15 -5969
rect 15 -4993 73 -4981
rect 15 -5969 27 -4993
rect 61 -5969 73 -4993
rect 15 -5981 73 -5969
<< ndiffc >>
rect -61 4993 -27 5969
rect 27 4993 61 5969
rect -61 3775 -27 4751
rect 27 3775 61 4751
rect -61 2557 -27 3533
rect 27 2557 61 3533
rect -61 1339 -27 2315
rect 27 1339 61 2315
rect -61 121 -27 1097
rect 27 121 61 1097
rect -61 -1097 -27 -121
rect 27 -1097 61 -121
rect -61 -2315 -27 -1339
rect 27 -2315 61 -1339
rect -61 -3533 -27 -2557
rect 27 -3533 61 -2557
rect -61 -4751 -27 -3775
rect 27 -4751 61 -3775
rect -61 -5969 -27 -4993
rect 27 -5969 61 -4993
<< psubdiff >>
rect -175 6121 -79 6155
rect 79 6121 175 6155
rect -175 6059 -141 6121
rect 141 6059 175 6121
rect -175 -6121 -141 -6059
rect 141 -6121 175 -6059
rect -175 -6155 -79 -6121
rect 79 -6155 175 -6121
<< psubdiffcont >>
rect -79 6121 79 6155
rect -175 -6059 -141 6059
rect 141 -6059 175 6059
rect -79 -6155 79 -6121
<< poly >>
rect -33 6053 33 6069
rect -33 6019 -17 6053
rect 17 6019 33 6053
rect -33 6003 33 6019
rect -15 5981 15 6003
rect -15 4959 15 4981
rect -33 4943 33 4959
rect -33 4909 -17 4943
rect 17 4909 33 4943
rect -33 4893 33 4909
rect -33 4835 33 4851
rect -33 4801 -17 4835
rect 17 4801 33 4835
rect -33 4785 33 4801
rect -15 4763 15 4785
rect -15 3741 15 3763
rect -33 3725 33 3741
rect -33 3691 -17 3725
rect 17 3691 33 3725
rect -33 3675 33 3691
rect -33 3617 33 3633
rect -33 3583 -17 3617
rect 17 3583 33 3617
rect -33 3567 33 3583
rect -15 3545 15 3567
rect -15 2523 15 2545
rect -33 2507 33 2523
rect -33 2473 -17 2507
rect 17 2473 33 2507
rect -33 2457 33 2473
rect -33 2399 33 2415
rect -33 2365 -17 2399
rect 17 2365 33 2399
rect -33 2349 33 2365
rect -15 2327 15 2349
rect -15 1305 15 1327
rect -33 1289 33 1305
rect -33 1255 -17 1289
rect 17 1255 33 1289
rect -33 1239 33 1255
rect -33 1181 33 1197
rect -33 1147 -17 1181
rect 17 1147 33 1181
rect -33 1131 33 1147
rect -15 1109 15 1131
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -1131 15 -1109
rect -33 -1147 33 -1131
rect -33 -1181 -17 -1147
rect 17 -1181 33 -1147
rect -33 -1197 33 -1181
rect -33 -1255 33 -1239
rect -33 -1289 -17 -1255
rect 17 -1289 33 -1255
rect -33 -1305 33 -1289
rect -15 -1327 15 -1305
rect -15 -2349 15 -2327
rect -33 -2365 33 -2349
rect -33 -2399 -17 -2365
rect 17 -2399 33 -2365
rect -33 -2415 33 -2399
rect -33 -2473 33 -2457
rect -33 -2507 -17 -2473
rect 17 -2507 33 -2473
rect -33 -2523 33 -2507
rect -15 -2545 15 -2523
rect -15 -3567 15 -3545
rect -33 -3583 33 -3567
rect -33 -3617 -17 -3583
rect 17 -3617 33 -3583
rect -33 -3633 33 -3617
rect -33 -3691 33 -3675
rect -33 -3725 -17 -3691
rect 17 -3725 33 -3691
rect -33 -3741 33 -3725
rect -15 -3763 15 -3741
rect -15 -4785 15 -4763
rect -33 -4801 33 -4785
rect -33 -4835 -17 -4801
rect 17 -4835 33 -4801
rect -33 -4851 33 -4835
rect -33 -4909 33 -4893
rect -33 -4943 -17 -4909
rect 17 -4943 33 -4909
rect -33 -4959 33 -4943
rect -15 -4981 15 -4959
rect -15 -6003 15 -5981
rect -33 -6019 33 -6003
rect -33 -6053 -17 -6019
rect 17 -6053 33 -6019
rect -33 -6069 33 -6053
<< polycont >>
rect -17 6019 17 6053
rect -17 4909 17 4943
rect -17 4801 17 4835
rect -17 3691 17 3725
rect -17 3583 17 3617
rect -17 2473 17 2507
rect -17 2365 17 2399
rect -17 1255 17 1289
rect -17 1147 17 1181
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -1181 17 -1147
rect -17 -1289 17 -1255
rect -17 -2399 17 -2365
rect -17 -2507 17 -2473
rect -17 -3617 17 -3583
rect -17 -3725 17 -3691
rect -17 -4835 17 -4801
rect -17 -4943 17 -4909
rect -17 -6053 17 -6019
<< locali >>
rect -175 6121 -79 6155
rect 79 6121 175 6155
rect -175 6059 -141 6121
rect 141 6059 175 6121
rect -33 6019 -17 6053
rect 17 6019 33 6053
rect -61 5969 -27 5985
rect -61 4977 -27 4993
rect 27 5969 61 5985
rect 27 4977 61 4993
rect -33 4909 -17 4943
rect 17 4909 33 4943
rect -33 4801 -17 4835
rect 17 4801 33 4835
rect -61 4751 -27 4767
rect -61 3759 -27 3775
rect 27 4751 61 4767
rect 27 3759 61 3775
rect -33 3691 -17 3725
rect 17 3691 33 3725
rect -33 3583 -17 3617
rect 17 3583 33 3617
rect -61 3533 -27 3549
rect -61 2541 -27 2557
rect 27 3533 61 3549
rect 27 2541 61 2557
rect -33 2473 -17 2507
rect 17 2473 33 2507
rect -33 2365 -17 2399
rect 17 2365 33 2399
rect -61 2315 -27 2331
rect -61 1323 -27 1339
rect 27 2315 61 2331
rect 27 1323 61 1339
rect -33 1255 -17 1289
rect 17 1255 33 1289
rect -33 1147 -17 1181
rect 17 1147 33 1181
rect -61 1097 -27 1113
rect -61 105 -27 121
rect 27 1097 61 1113
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -1113 -27 -1097
rect 27 -121 61 -105
rect 27 -1113 61 -1097
rect -33 -1181 -17 -1147
rect 17 -1181 33 -1147
rect -33 -1289 -17 -1255
rect 17 -1289 33 -1255
rect -61 -1339 -27 -1323
rect -61 -2331 -27 -2315
rect 27 -1339 61 -1323
rect 27 -2331 61 -2315
rect -33 -2399 -17 -2365
rect 17 -2399 33 -2365
rect -33 -2507 -17 -2473
rect 17 -2507 33 -2473
rect -61 -2557 -27 -2541
rect -61 -3549 -27 -3533
rect 27 -2557 61 -2541
rect 27 -3549 61 -3533
rect -33 -3617 -17 -3583
rect 17 -3617 33 -3583
rect -33 -3725 -17 -3691
rect 17 -3725 33 -3691
rect -61 -3775 -27 -3759
rect -61 -4767 -27 -4751
rect 27 -3775 61 -3759
rect 27 -4767 61 -4751
rect -33 -4835 -17 -4801
rect 17 -4835 33 -4801
rect -33 -4943 -17 -4909
rect 17 -4943 33 -4909
rect -61 -4993 -27 -4977
rect -61 -5985 -27 -5969
rect 27 -4993 61 -4977
rect 27 -5985 61 -5969
rect -33 -6053 -17 -6019
rect 17 -6053 33 -6019
rect -175 -6121 -141 -6059
rect 141 -6121 175 -6059
rect -175 -6155 -79 -6121
rect 79 -6155 175 -6121
<< viali >>
rect -17 6019 17 6053
rect -61 4993 -27 5969
rect 27 4993 61 5969
rect -17 4909 17 4943
rect -17 4801 17 4835
rect -61 3775 -27 4751
rect 27 3775 61 4751
rect -17 3691 17 3725
rect -17 3583 17 3617
rect -61 2557 -27 3533
rect 27 2557 61 3533
rect -17 2473 17 2507
rect -17 2365 17 2399
rect -61 1339 -27 2315
rect 27 1339 61 2315
rect -17 1255 17 1289
rect -17 1147 17 1181
rect -61 121 -27 1097
rect 27 121 61 1097
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -1097 -27 -121
rect 27 -1097 61 -121
rect -17 -1181 17 -1147
rect -17 -1289 17 -1255
rect -61 -2315 -27 -1339
rect 27 -2315 61 -1339
rect -17 -2399 17 -2365
rect -17 -2507 17 -2473
rect -61 -3533 -27 -2557
rect 27 -3533 61 -2557
rect -17 -3617 17 -3583
rect -17 -3725 17 -3691
rect -61 -4751 -27 -3775
rect 27 -4751 61 -3775
rect -17 -4835 17 -4801
rect -17 -4943 17 -4909
rect -61 -5969 -27 -4993
rect 27 -5969 61 -4993
rect -17 -6053 17 -6019
<< metal1 >>
rect -29 6053 29 6059
rect -29 6019 -17 6053
rect 17 6019 29 6053
rect -29 6013 29 6019
rect -67 5969 -21 5981
rect -67 4993 -61 5969
rect -27 4993 -21 5969
rect -67 4981 -21 4993
rect 21 5969 67 5981
rect 21 4993 27 5969
rect 61 4993 67 5969
rect 21 4981 67 4993
rect -29 4943 29 4949
rect -29 4909 -17 4943
rect 17 4909 29 4943
rect -29 4903 29 4909
rect -29 4835 29 4841
rect -29 4801 -17 4835
rect 17 4801 29 4835
rect -29 4795 29 4801
rect -67 4751 -21 4763
rect -67 3775 -61 4751
rect -27 3775 -21 4751
rect -67 3763 -21 3775
rect 21 4751 67 4763
rect 21 3775 27 4751
rect 61 3775 67 4751
rect 21 3763 67 3775
rect -29 3725 29 3731
rect -29 3691 -17 3725
rect 17 3691 29 3725
rect -29 3685 29 3691
rect -29 3617 29 3623
rect -29 3583 -17 3617
rect 17 3583 29 3617
rect -29 3577 29 3583
rect -67 3533 -21 3545
rect -67 2557 -61 3533
rect -27 2557 -21 3533
rect -67 2545 -21 2557
rect 21 3533 67 3545
rect 21 2557 27 3533
rect 61 2557 67 3533
rect 21 2545 67 2557
rect -29 2507 29 2513
rect -29 2473 -17 2507
rect 17 2473 29 2507
rect -29 2467 29 2473
rect -29 2399 29 2405
rect -29 2365 -17 2399
rect 17 2365 29 2399
rect -29 2359 29 2365
rect -67 2315 -21 2327
rect -67 1339 -61 2315
rect -27 1339 -21 2315
rect -67 1327 -21 1339
rect 21 2315 67 2327
rect 21 1339 27 2315
rect 61 1339 67 2315
rect 21 1327 67 1339
rect -29 1289 29 1295
rect -29 1255 -17 1289
rect 17 1255 29 1289
rect -29 1249 29 1255
rect -29 1181 29 1187
rect -29 1147 -17 1181
rect 17 1147 29 1181
rect -29 1141 29 1147
rect -67 1097 -21 1109
rect -67 121 -61 1097
rect -27 121 -21 1097
rect -67 109 -21 121
rect 21 1097 67 1109
rect 21 121 27 1097
rect 61 121 67 1097
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -1097 -61 -121
rect -27 -1097 -21 -121
rect -67 -1109 -21 -1097
rect 21 -121 67 -109
rect 21 -1097 27 -121
rect 61 -1097 67 -121
rect 21 -1109 67 -1097
rect -29 -1147 29 -1141
rect -29 -1181 -17 -1147
rect 17 -1181 29 -1147
rect -29 -1187 29 -1181
rect -29 -1255 29 -1249
rect -29 -1289 -17 -1255
rect 17 -1289 29 -1255
rect -29 -1295 29 -1289
rect -67 -1339 -21 -1327
rect -67 -2315 -61 -1339
rect -27 -2315 -21 -1339
rect -67 -2327 -21 -2315
rect 21 -1339 67 -1327
rect 21 -2315 27 -1339
rect 61 -2315 67 -1339
rect 21 -2327 67 -2315
rect -29 -2365 29 -2359
rect -29 -2399 -17 -2365
rect 17 -2399 29 -2365
rect -29 -2405 29 -2399
rect -29 -2473 29 -2467
rect -29 -2507 -17 -2473
rect 17 -2507 29 -2473
rect -29 -2513 29 -2507
rect -67 -2557 -21 -2545
rect -67 -3533 -61 -2557
rect -27 -3533 -21 -2557
rect -67 -3545 -21 -3533
rect 21 -2557 67 -2545
rect 21 -3533 27 -2557
rect 61 -3533 67 -2557
rect 21 -3545 67 -3533
rect -29 -3583 29 -3577
rect -29 -3617 -17 -3583
rect 17 -3617 29 -3583
rect -29 -3623 29 -3617
rect -29 -3691 29 -3685
rect -29 -3725 -17 -3691
rect 17 -3725 29 -3691
rect -29 -3731 29 -3725
rect -67 -3775 -21 -3763
rect -67 -4751 -61 -3775
rect -27 -4751 -21 -3775
rect -67 -4763 -21 -4751
rect 21 -3775 67 -3763
rect 21 -4751 27 -3775
rect 61 -4751 67 -3775
rect 21 -4763 67 -4751
rect -29 -4801 29 -4795
rect -29 -4835 -17 -4801
rect 17 -4835 29 -4801
rect -29 -4841 29 -4835
rect -29 -4909 29 -4903
rect -29 -4943 -17 -4909
rect 17 -4943 29 -4909
rect -29 -4949 29 -4943
rect -67 -4993 -21 -4981
rect -67 -5969 -61 -4993
rect -27 -5969 -21 -4993
rect -67 -5981 -21 -5969
rect 21 -4993 67 -4981
rect 21 -5969 27 -4993
rect 61 -5969 67 -4993
rect 21 -5981 67 -5969
rect -29 -6019 29 -6013
rect -29 -6053 -17 -6019
rect 17 -6053 29 -6019
rect -29 -6059 29 -6053
<< properties >>
string FIXED_BBOX -158 -6138 158 6138
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
