magic
tech sky130A
magscale 1 2
timestamp 1666052912
<< metal4 >>
rect -10447 959 -3749 1000
rect -10447 481 -4005 959
rect -3769 481 -3749 959
rect -10447 440 -3749 481
rect -3349 959 3349 1000
rect -3349 481 3093 959
rect 3329 481 3349 959
rect -3349 440 3349 481
rect 3749 959 10447 1000
rect 3749 481 10191 959
rect 10427 481 10447 959
rect 3749 440 10447 481
rect -10447 239 -3749 280
rect -10447 -239 -4005 239
rect -3769 -239 -3749 239
rect -10447 -280 -3749 -239
rect -3349 239 3349 280
rect -3349 -239 3093 239
rect 3329 -239 3349 239
rect -3349 -280 3349 -239
rect 3749 239 10447 280
rect 3749 -239 10191 239
rect 10427 -239 10447 239
rect 3749 -280 10447 -239
rect -10447 -481 -3749 -440
rect -10447 -959 -4005 -481
rect -3769 -959 -3749 -481
rect -10447 -1000 -3749 -959
rect -3349 -481 3349 -440
rect -3349 -959 3093 -481
rect 3329 -959 3349 -481
rect -3349 -1000 3349 -959
rect 3749 -481 10447 -440
rect 3749 -959 10191 -481
rect 10427 -959 10447 -481
rect 3749 -1000 10447 -959
<< via4 >>
rect -4005 481 -3769 959
rect 3093 481 3329 959
rect 10191 481 10427 959
rect -4005 -239 -3769 239
rect 3093 -239 3329 239
rect 10191 -239 10427 239
rect -4005 -959 -3769 -481
rect 3093 -959 3329 -481
rect 10191 -959 10427 -481
<< mimcap2 >>
rect -10367 880 -4367 920
rect -10367 560 -10327 880
rect -4407 560 -4367 880
rect -10367 520 -4367 560
rect -3269 880 2731 920
rect -3269 560 -3229 880
rect 2691 560 2731 880
rect -3269 520 2731 560
rect 3829 880 9829 920
rect 3829 560 3869 880
rect 9789 560 9829 880
rect 3829 520 9829 560
rect -10367 160 -4367 200
rect -10367 -160 -10327 160
rect -4407 -160 -4367 160
rect -10367 -200 -4367 -160
rect -3269 160 2731 200
rect -3269 -160 -3229 160
rect 2691 -160 2731 160
rect -3269 -200 2731 -160
rect 3829 160 9829 200
rect 3829 -160 3869 160
rect 9789 -160 9829 160
rect 3829 -200 9829 -160
rect -10367 -560 -4367 -520
rect -10367 -880 -10327 -560
rect -4407 -880 -4367 -560
rect -10367 -920 -4367 -880
rect -3269 -560 2731 -520
rect -3269 -880 -3229 -560
rect 2691 -880 2731 -560
rect -3269 -920 2731 -880
rect 3829 -560 9829 -520
rect 3829 -880 3869 -560
rect 9789 -880 9829 -560
rect 3829 -920 9829 -880
<< mimcap2contact >>
rect -10327 560 -4407 880
rect -3229 560 2691 880
rect 3869 560 9789 880
rect -10327 -160 -4407 160
rect -3229 -160 2691 160
rect 3869 -160 9789 160
rect -10327 -880 -4407 -560
rect -3229 -880 2691 -560
rect 3869 -880 9789 -560
<< metal5 >>
rect -7527 904 -7207 1080
rect -4047 959 -3727 1080
rect -10351 880 -4383 904
rect -10351 560 -10327 880
rect -4407 560 -4383 880
rect -10351 536 -4383 560
rect -7527 184 -7207 536
rect -4047 481 -4005 959
rect -3769 481 -3727 959
rect -429 904 -109 1080
rect 3051 959 3371 1080
rect -3253 880 2715 904
rect -3253 560 -3229 880
rect 2691 560 2715 880
rect -3253 536 2715 560
rect -4047 239 -3727 481
rect -10351 160 -4383 184
rect -10351 -160 -10327 160
rect -4407 -160 -4383 160
rect -10351 -184 -4383 -160
rect -7527 -536 -7207 -184
rect -4047 -239 -4005 239
rect -3769 -239 -3727 239
rect -429 184 -109 536
rect 3051 481 3093 959
rect 3329 481 3371 959
rect 6669 904 6989 1080
rect 10149 959 10469 1080
rect 3845 880 9813 904
rect 3845 560 3869 880
rect 9789 560 9813 880
rect 3845 536 9813 560
rect 3051 239 3371 481
rect -3253 160 2715 184
rect -3253 -160 -3229 160
rect 2691 -160 2715 160
rect -3253 -184 2715 -160
rect -4047 -481 -3727 -239
rect -10351 -560 -4383 -536
rect -10351 -880 -10327 -560
rect -4407 -880 -4383 -560
rect -10351 -904 -4383 -880
rect -7527 -1080 -7207 -904
rect -4047 -959 -4005 -481
rect -3769 -959 -3727 -481
rect -429 -536 -109 -184
rect 3051 -239 3093 239
rect 3329 -239 3371 239
rect 6669 184 6989 536
rect 10149 481 10191 959
rect 10427 481 10469 959
rect 10149 239 10469 481
rect 3845 160 9813 184
rect 3845 -160 3869 160
rect 9789 -160 9813 160
rect 3845 -184 9813 -160
rect 3051 -481 3371 -239
rect -3253 -560 2715 -536
rect -3253 -880 -3229 -560
rect 2691 -880 2715 -560
rect -3253 -904 2715 -880
rect -4047 -1080 -3727 -959
rect -429 -1080 -109 -904
rect 3051 -959 3093 -481
rect 3329 -959 3371 -481
rect 6669 -536 6989 -184
rect 10149 -239 10191 239
rect 10427 -239 10469 239
rect 10149 -481 10469 -239
rect 3845 -560 9813 -536
rect 3845 -880 3869 -560
rect 9789 -880 9813 -560
rect 3845 -904 9813 -880
rect 3051 -1080 3371 -959
rect 6669 -1080 6989 -904
rect 10149 -959 10191 -481
rect 10427 -959 10469 -481
rect 10149 -1080 10469 -959
<< properties >>
string FIXED_BBOX 3749 440 9909 1000
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30.0 l 2.00 val 132.16 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
