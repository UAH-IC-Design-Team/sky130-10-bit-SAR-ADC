magic
tech sky130A
timestamp 1666625366
<< metal1 >>
rect 0 0 10000 10000
<< end >>
