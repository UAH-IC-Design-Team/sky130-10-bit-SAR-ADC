magic
tech sky130A
magscale 1 2
timestamp 1666649035
<< metal3 >>
rect -1150 10272 1149 10300
rect -1150 8128 1065 10272
rect 1129 8128 1149 10272
rect -1150 8100 1149 8128
rect -1150 7972 1149 8000
rect -1150 5828 1065 7972
rect 1129 5828 1149 7972
rect -1150 5800 1149 5828
rect -1150 5672 1149 5700
rect -1150 3528 1065 5672
rect 1129 3528 1149 5672
rect -1150 3500 1149 3528
rect -1150 3372 1149 3400
rect -1150 1228 1065 3372
rect 1129 2179 1149 3372
rect 1129 1228 2305 2179
rect -1150 1200 2305 1228
rect 6 1100 2305 1200
rect -1150 1072 2305 1100
rect -1150 -1072 1065 1072
rect 1129 -21 2305 1072
rect 1129 -1072 1149 -21
rect -1150 -1100 1149 -1072
rect -1150 -1228 1149 -1200
rect -1150 -3372 1065 -1228
rect 1129 -3372 1149 -1228
rect -1150 -3400 1149 -3372
rect -1150 -3528 1149 -3500
rect -1150 -5672 1065 -3528
rect 1129 -5672 1149 -3528
rect -1150 -5700 1149 -5672
rect -1150 -5828 1149 -5800
rect -1150 -7972 1065 -5828
rect 1129 -7972 1149 -5828
rect -1150 -8000 1149 -7972
rect -1150 -8128 1149 -8100
rect -1150 -10272 1065 -8128
rect 1129 -10272 1149 -8128
rect -1150 -10300 1149 -10272
<< via3 >>
rect 1065 8128 1129 10272
rect 1065 5828 1129 7972
rect 1065 3528 1129 5672
rect 1065 1228 1129 3372
rect 1065 -1072 1129 1072
rect 1065 -3372 1129 -1228
rect 1065 -5672 1129 -3528
rect 1065 -7972 1129 -5828
rect 1065 -10272 1129 -8128
<< mimcap >>
rect -1050 10160 950 10200
rect -1050 8240 -1010 10160
rect 910 8240 950 10160
rect -1050 8200 950 8240
rect -1050 7860 950 7900
rect -1050 5940 -1010 7860
rect 910 5940 950 7860
rect -1050 5900 950 5940
rect -1050 5560 950 5600
rect -1050 3640 -1010 5560
rect 910 3640 950 5560
rect -1050 3600 950 3640
rect -1050 3260 950 3300
rect -1050 1340 -1010 3260
rect 910 1340 950 3260
rect -1050 1300 950 1340
rect -1050 960 950 1000
rect -1050 -960 -1010 960
rect 910 -960 950 960
rect -1050 -1000 950 -960
rect -1050 -1340 950 -1300
rect -1050 -3260 -1010 -1340
rect 910 -3260 950 -1340
rect -1050 -3300 950 -3260
rect -1050 -3640 950 -3600
rect -1050 -5560 -1010 -3640
rect 910 -5560 950 -3640
rect -1050 -5600 950 -5560
rect -1050 -5940 950 -5900
rect -1050 -7860 -1010 -5940
rect 910 -7860 950 -5940
rect -1050 -7900 950 -7860
rect -1050 -8240 950 -8200
rect -1050 -10160 -1010 -8240
rect 910 -10160 950 -8240
rect -1050 -10200 950 -10160
<< mimcapcontact >>
rect -1010 8240 910 10160
rect -1010 5940 910 7860
rect -1010 3640 910 5560
rect -1010 1340 910 3260
rect -1010 -960 910 960
rect -1010 -3260 910 -1340
rect -1010 -5560 910 -3640
rect -1010 -7860 910 -5940
rect -1010 -10160 910 -8240
<< metal4 >>
rect -102 10161 2 10350
rect 1018 10288 1122 10350
rect 1018 10272 1145 10288
rect -1011 10160 911 10161
rect -1011 8240 -1010 10160
rect 910 8240 911 10160
rect -1011 8239 911 8240
rect -102 7861 2 8239
rect 1018 8128 1065 10272
rect 1129 8128 1145 10272
rect 1018 8112 1145 8128
rect 1018 7988 1122 8112
rect 1018 7972 1145 7988
rect -1011 7860 911 7861
rect -1011 5940 -1010 7860
rect 910 5940 911 7860
rect -1011 5939 911 5940
rect -102 5561 2 5939
rect 1018 5828 1065 7972
rect 1129 5828 1145 7972
rect 1018 5812 1145 5828
rect 1018 5688 1122 5812
rect 1018 5672 1145 5688
rect -1011 5560 911 5561
rect -1011 3640 -1010 5560
rect 910 3640 911 5560
rect -1011 3639 911 3640
rect -102 3261 2 3639
rect 1018 3528 1065 5672
rect 1129 3528 1145 5672
rect 1018 3512 1145 3528
rect 1018 3388 1122 3512
rect 1018 3372 1145 3388
rect -1011 3260 911 3261
rect -1011 1340 -1010 3260
rect 910 1340 911 3260
rect -1011 1339 911 1340
rect -102 961 2 1339
rect 1018 1228 1065 3372
rect 1129 1228 1145 3372
rect 1018 1212 1145 1228
rect 1018 1088 1122 1212
rect 1018 1072 1145 1088
rect -1011 960 911 961
rect -1011 -960 -1010 960
rect 910 -960 911 960
rect -1011 -961 911 -960
rect -102 -1339 2 -961
rect 1018 -1072 1065 1072
rect 1129 -1072 1145 1072
rect 1018 -1088 1145 -1072
rect 1018 -1212 1122 -1088
rect 1018 -1228 1145 -1212
rect -1011 -1340 911 -1339
rect -1011 -3260 -1010 -1340
rect 910 -3260 911 -1340
rect -1011 -3261 911 -3260
rect -102 -3639 2 -3261
rect 1018 -3372 1065 -1228
rect 1129 -3372 1145 -1228
rect 1018 -3388 1145 -3372
rect 1018 -3512 1122 -3388
rect 1018 -3528 1145 -3512
rect -1011 -3640 911 -3639
rect -1011 -5560 -1010 -3640
rect 910 -5560 911 -3640
rect -1011 -5561 911 -5560
rect -102 -5939 2 -5561
rect 1018 -5672 1065 -3528
rect 1129 -5672 1145 -3528
rect 1018 -5688 1145 -5672
rect 1018 -5812 1122 -5688
rect 1018 -5828 1145 -5812
rect -1011 -5940 911 -5939
rect -1011 -7860 -1010 -5940
rect 910 -7860 911 -5940
rect -1011 -7861 911 -7860
rect -102 -8239 2 -7861
rect 1018 -7972 1065 -5828
rect 1129 -7972 1145 -5828
rect 1018 -7988 1145 -7972
rect 1018 -8112 1122 -7988
rect 1018 -8128 1145 -8112
rect -1011 -8240 911 -8239
rect -1011 -10160 -1010 -8240
rect 910 -10160 911 -8240
rect -1011 -10161 911 -10160
rect -102 -10350 2 -10161
rect 1018 -10272 1065 -8128
rect 1129 -10272 1145 -8128
rect 1018 -10288 1145 -10272
rect 1018 -10350 1122 -10288
<< properties >>
string FIXED_BBOX -1150 8100 1050 10300
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 9 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
