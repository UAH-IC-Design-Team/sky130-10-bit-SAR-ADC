magic
tech sky130A
magscale 1 2
timestamp 1668286849
<< metal1 >>
rect 138240 31400 160990 31460
rect 161220 31400 161240 31460
rect 138140 28490 138200 28500
rect 138140 25360 138200 28290
rect 133700 25300 138200 25360
rect 138240 25260 138300 31400
rect 133700 25200 138300 25260
rect 138340 31300 159690 31360
rect 159930 31300 159950 31360
rect 138340 25160 138400 31300
rect 133700 25100 138400 25160
rect 138440 31200 158410 31260
rect 158650 31200 158660 31260
rect 138440 25060 138500 31200
rect 133700 25000 138500 25060
rect 138540 31100 157130 31160
rect 157360 31100 157370 31160
rect 138540 24960 138600 31100
rect 133700 24900 138600 24960
rect 138640 31000 155830 31060
rect 156070 31000 156080 31060
rect 138640 24860 138700 31000
rect 133700 24800 138700 24860
rect 138740 30900 154550 30960
rect 154780 30900 154800 30960
rect 138740 24760 138800 30900
rect 133700 24700 138800 24760
rect 138840 30800 153280 30860
rect 153490 30800 153510 30860
rect 138840 24660 138900 30800
rect 133700 24600 138900 24660
rect 138940 30700 151990 30760
rect 152210 30700 152220 30760
rect 138940 24560 139000 30700
rect 133700 24500 139000 24560
rect 139040 30600 150690 30660
rect 150920 30600 150930 30660
rect 139040 24460 139100 30600
rect 133700 24400 139100 24460
rect 139140 30500 149390 30560
rect 149630 30500 149640 30560
rect 139140 24360 139200 30500
rect 133700 24300 139200 24360
rect 139240 30400 148130 30460
rect 148340 30400 148400 30460
rect 139240 24260 139300 30400
rect 133700 24200 139300 24260
rect 139340 30300 146870 30360
rect 147070 30300 147080 30360
rect 139340 24160 139400 30300
rect 133700 24100 139400 24160
rect 139440 30200 145590 30260
rect 145790 30200 145800 30260
rect 139440 24060 139500 30200
rect 133700 24000 139500 24060
rect 139540 30100 144290 30160
rect 144490 30100 144500 30160
rect 139540 23960 139600 30100
rect 133700 23900 139600 23960
rect 139640 30000 142990 30060
rect 143190 30000 143200 30060
rect 139640 23860 139700 30000
rect 133700 23800 139700 23860
rect 139740 29900 141710 29960
rect 141910 29900 141920 29960
rect 139740 23760 139800 29900
rect 133700 23700 139800 23760
rect 139840 29800 140430 29860
rect 140630 29800 140640 29860
rect 139840 23660 139900 29800
rect 140000 28480 140500 28500
rect 140000 28380 140020 28480
rect 140480 28380 140500 28480
rect 140060 28360 140500 28380
rect 133700 23600 139900 23660
rect 137400 23390 137600 23400
rect 137400 23010 137410 23390
rect 137590 23010 137600 23390
rect 137400 23000 137600 23010
rect 1490 19490 1710 19860
rect 1490 17690 1710 18060
rect 137400 14610 137590 14620
rect 137400 14330 137410 14610
rect 137580 14330 137590 14610
rect 137400 14320 137590 14330
rect 138840 14240 138860 14380
rect 138940 14240 138960 14380
rect 138840 14220 138960 14240
rect 133700 13740 139900 13800
rect 133700 13640 139800 13700
rect 133700 13540 139700 13600
rect 133700 13440 139600 13500
rect 133700 13340 139500 13400
rect 133700 13240 139400 13300
rect 133700 13140 139300 13200
rect 133700 13040 139200 13100
rect 133700 12940 139100 13000
rect 133700 12840 139000 12900
rect 133700 12740 138900 12800
rect 133700 12640 138800 12700
rect 133700 12540 138700 12600
rect 133700 12440 138600 12500
rect 133700 12340 138500 12400
rect 133700 12240 138400 12300
rect 133700 12140 138300 12200
rect 138240 6000 138300 12140
rect 138340 6100 138400 12240
rect 138440 6200 138500 12340
rect 138540 6300 138600 12440
rect 138640 6400 138700 12540
rect 138740 6500 138800 12640
rect 138840 6600 138900 12740
rect 138940 6700 139000 12840
rect 139040 6800 139100 12940
rect 139140 6900 139200 13040
rect 139240 7000 139300 13140
rect 139340 7100 139400 13240
rect 139440 7200 139500 13340
rect 139540 7300 139600 13440
rect 139640 7400 139700 13540
rect 139740 7500 139800 13640
rect 139840 7600 139900 13740
rect 139840 7540 140350 7600
rect 140610 7540 140620 7600
rect 139740 7440 141610 7500
rect 141870 7440 141900 7500
rect 139640 7340 142910 7400
rect 143190 7340 143220 7400
rect 139540 7240 144230 7300
rect 144480 7240 144520 7300
rect 139440 7140 145470 7200
rect 145770 7140 145820 7200
rect 139340 7040 146770 7100
rect 147060 7040 147100 7100
rect 139240 6940 148050 7000
rect 148340 6940 148400 7000
rect 139140 6840 149350 6900
rect 149630 6840 149660 6900
rect 139040 6740 150610 6800
rect 150920 6740 150960 6800
rect 138940 6640 151930 6700
rect 152210 6640 152260 6700
rect 138840 6540 153210 6600
rect 153490 6540 153560 6600
rect 138740 6440 154490 6500
rect 154780 6440 154820 6500
rect 138640 6340 155770 6400
rect 156060 6340 156100 6400
rect 138540 6240 157050 6300
rect 157360 6240 157400 6300
rect 138440 6140 158350 6200
rect 158650 6140 158680 6200
rect 138340 6040 159630 6100
rect 159930 6040 159960 6100
rect 138240 5940 160930 6000
rect 161220 5940 161260 6000
<< via1 >>
rect 160990 31400 161220 31460
rect 138140 28290 138200 28490
rect 159690 31300 159930 31360
rect 158410 31200 158650 31260
rect 157130 31100 157360 31160
rect 155830 31000 156070 31060
rect 154550 30900 154780 30960
rect 153280 30800 153490 30860
rect 151990 30700 152210 30760
rect 150690 30600 150920 30660
rect 149390 30500 149630 30560
rect 148130 30400 148340 30460
rect 146870 30300 147070 30360
rect 145590 30200 145790 30260
rect 144290 30100 144490 30160
rect 142990 30000 143190 30060
rect 141710 29900 141910 29960
rect 140430 29800 140630 29860
rect 140020 28380 140480 28480
rect 137410 23010 137590 23390
rect 137410 14330 137580 14610
rect 138860 14240 138940 14440
rect 140350 7540 140610 7600
rect 141610 7440 141870 7500
rect 142910 7340 143190 7400
rect 144230 7240 144480 7300
rect 145470 7140 145770 7200
rect 146770 7040 147060 7100
rect 148050 6940 148340 7000
rect 149350 6840 149630 6900
rect 150610 6740 150920 6800
rect 151930 6640 152210 6700
rect 153210 6540 153490 6600
rect 154490 6440 154780 6500
rect 155770 6340 156060 6400
rect 157050 6240 157360 6300
rect 158350 6140 158650 6200
rect 159630 6040 159930 6100
rect 160930 5940 161220 6000
<< metal2 >>
rect 161178 31460 161234 31465
rect 160980 31400 160990 31460
rect 161220 31400 161234 31460
rect 159890 31360 159946 31365
rect 159680 31300 159690 31360
rect 159930 31300 159946 31360
rect 158602 31260 158658 31265
rect 158400 31200 158410 31260
rect 158650 31200 158658 31260
rect 157314 31160 157370 31165
rect 157120 31100 157130 31160
rect 157360 31100 157370 31160
rect 156026 31060 156082 31065
rect 155820 31000 155830 31060
rect 156070 31000 156082 31060
rect 154738 30960 154794 30965
rect 154540 30900 154550 30960
rect 154780 30900 154794 30960
rect 153450 30860 153506 30865
rect 153260 30800 153280 30860
rect 153490 30800 153506 30860
rect 152162 30760 152218 30765
rect 151980 30700 151990 30760
rect 152210 30700 152218 30760
rect 150874 30660 150930 30665
rect 150680 30600 150690 30660
rect 150920 30600 150930 30660
rect 149380 30500 149390 30560
rect 148120 30400 148130 30460
rect 146860 30300 146870 30360
rect 147070 30300 147080 30360
rect 145580 30200 145590 30260
rect 145790 30200 145800 30260
rect 144280 30100 144290 30160
rect 144490 30100 144500 30160
rect 142980 30000 142990 30060
rect 143190 30000 143200 30060
rect 141700 29900 141710 29960
rect 141910 29900 141920 29960
rect 150874 29865 150930 30600
rect 152162 29965 152218 30700
rect 153450 30065 153506 30800
rect 154738 30165 154794 30900
rect 140420 29800 140430 29860
rect 140630 29800 140640 29860
rect 156026 29845 156082 31000
rect 157314 30365 157370 31100
rect 158602 30465 158658 31200
rect 159890 30565 159946 31300
rect 161178 30565 161234 31400
rect 138140 28490 140500 28500
rect 138200 28480 140500 28490
rect 138200 28380 140020 28480
rect 140480 28380 140500 28480
rect 138200 28360 140500 28380
rect 138140 28280 138200 28290
rect 137400 23390 137600 23400
rect 137400 23010 137410 23390
rect 137590 23010 137600 23390
rect 137400 23000 137600 23010
rect 137400 14610 137590 14620
rect 137400 14330 137410 14610
rect 137580 14330 137590 14610
rect 137400 14320 137590 14330
rect 138820 14440 138980 14480
rect 138820 14240 138860 14440
rect 138940 14240 138980 14440
rect 138820 8780 138980 14240
rect 138820 8760 140540 8780
rect 138820 8660 140010 8760
rect 140530 8660 140540 8760
rect 138820 8640 140540 8660
rect 140340 7540 140350 7600
rect 140610 7540 140620 7600
rect 141600 7440 141610 7500
rect 141870 7440 141880 7500
rect 142900 7340 142910 7400
rect 144220 7240 144230 7300
rect 144480 7240 144500 7300
rect 145460 7140 145470 7200
rect 146760 7040 146770 7100
rect 148040 6940 148050 7000
rect 149340 6840 149350 6900
rect 150600 6740 150610 6800
rect 151920 6640 151930 6700
rect 153450 6600 153506 7340
rect 153200 6540 153210 6600
rect 153490 6540 153506 6600
rect 154738 6500 154794 7240
rect 154480 6440 154490 6500
rect 154780 6440 154794 6500
rect 156026 6400 156082 7140
rect 155760 6340 155770 6400
rect 156060 6340 156082 6400
rect 157314 6300 157370 7040
rect 157040 6240 157050 6300
rect 157360 6240 157370 6300
rect 158602 6200 158658 6940
rect 158340 6140 158350 6200
rect 158650 6140 158658 6200
rect 159890 6100 159946 6840
rect 159620 6040 159630 6100
rect 159930 6040 159946 6100
rect 161178 6000 161234 6740
rect 160920 5940 160930 6000
rect 161220 5940 161234 6000
<< via2 >>
rect 140020 28380 140480 28480
rect 137410 23010 137590 23390
rect 137410 14330 137580 14610
rect 140010 8660 140530 8760
<< metal3 >>
rect 161061 29184 161861 29304
rect 161061 27416 161861 27536
rect 134400 25980 136000 26000
rect 134400 25620 135220 25980
rect 135980 25620 136000 25980
rect 161061 25648 161861 25768
rect 134400 25600 136000 25620
rect 161061 23880 161861 24000
rect 137400 23400 140200 23600
rect 137400 23390 137600 23400
rect 137400 23010 137410 23390
rect 137590 23010 137600 23390
rect 137400 23000 137600 23010
rect 140000 20600 140200 23400
rect 161061 22112 161861 22232
rect 161061 20344 161861 20464
rect 161061 18576 161861 18696
rect 161061 16808 161861 16928
rect 137400 14610 137590 14620
rect 137400 14330 137410 14610
rect 137580 14330 137590 14610
rect 137400 13800 137590 14330
rect 140000 13800 140200 16600
rect 161061 15040 161861 15160
rect 137400 13600 140200 13800
rect 161061 13272 161861 13392
rect 134400 11660 136000 11700
rect 134400 11340 135240 11660
rect 135960 11340 136000 11660
rect 161061 11504 161861 11624
rect 134400 11300 136000 11340
rect 161284 9736 161861 9856
rect 161061 7968 161861 8088
<< via3 >>
rect 135220 25620 135980 25980
rect 135240 11340 135960 11660
<< metal4 >>
rect 140600 27360 141000 27400
rect 140600 27040 140640 27360
rect 140960 27040 141000 27360
rect 140600 26000 141000 27040
rect 135200 25980 141000 26000
rect 135200 25620 135220 25980
rect 135980 25620 141000 25980
rect 135200 25600 141000 25620
rect 135200 11660 141000 11700
rect 135200 11340 135240 11660
rect 135960 11340 141000 11660
rect 135200 11300 141000 11340
rect 140600 10560 141000 11300
rect 140600 10240 140640 10560
rect 140960 10240 141000 10560
rect 140600 10200 141000 10240
<< via4 >>
rect 140640 27040 140960 27360
rect 145840 27040 146160 27360
rect 150740 27040 151060 27360
rect 155640 27040 155960 27360
rect 160540 27040 160860 27360
rect 133640 25640 134360 25960
rect 143400 25640 143700 25960
rect 148300 25640 148600 25960
rect 153200 25640 153500 25960
rect 158100 25640 158400 25960
rect 133640 11340 134360 11660
rect 143400 11340 143700 11660
rect 148300 11340 148600 11660
rect 153200 11340 153500 11660
rect 158100 11340 158400 11660
rect 140640 10240 140960 10560
rect 145840 10240 146160 10560
rect 150740 10240 151060 10560
rect 155640 10240 155960 10560
rect 160540 10240 160860 10560
<< metal5 >>
rect 140600 27360 161000 27400
rect 140600 27040 140640 27360
rect 140960 27040 145840 27360
rect 146160 27040 150740 27360
rect 151060 27040 155640 27360
rect 155960 27040 160540 27360
rect 160860 27040 161000 27360
rect 140600 27000 161000 27040
rect 133600 25960 161000 26000
rect 133600 25640 133640 25960
rect 134360 25640 143400 25960
rect 143700 25640 148300 25960
rect 148600 25640 153200 25960
rect 153500 25640 158100 25960
rect 158400 25640 161000 25960
rect 133600 25600 161000 25640
rect 133600 11660 161000 11700
rect 133600 11340 133640 11660
rect 134360 11340 143400 11660
rect 143700 11340 148300 11660
rect 148600 11340 153200 11660
rect 153500 11340 158100 11660
rect 158400 11340 161000 11660
rect 133600 11300 161000 11340
rect 140600 10560 161000 10600
rect 140600 10240 140640 10560
rect 140960 10240 145840 10560
rect 146160 10240 150740 10560
rect 151060 10240 155640 10560
rect 155960 10240 160540 10560
rect 160860 10240 161000 10560
rect 140600 10200 161000 10240
use all_analog  all_analog_0 components
timestamp 1668283997
transform 1 0 5843800 0 1 6591400
box -5842300 -6591400 -5704620 -6554100
use controller  controller_0 components
timestamp 1668286574
transform 1 0 140000 0 1 6600
box 0 0 21861 24005
<< labels >>
rlabel metal5 158400 11300 161000 11700 1 VDD
port 1 n
rlabel metal1 1490 19490 1710 19860 1 V_in_p
port 2 n
rlabel metal3 161061 25648 161861 25768 1 Done
port 3 n
rlabel metal5 160860 10200 161000 10600 1 VSS
port 4 n
rlabel metal1 1490 17690 1710 18060 1 V_in_n
port 5 n
rlabel metal3 161061 27416 161861 27536 1 Clk
port 6 n
rlabel metal3 161061 7968 161861 8088 1 Bit10
port 7 n
rlabel metal3 161284 9736 161861 9856 1 Bit9
port 8 n
rlabel metal3 161061 11504 161861 11624 1 Bit8
port 9 n
rlabel metal3 161061 13272 161861 13392 1 Bit7
port 10 n
rlabel metal3 161061 15040 161861 15160 1 Bit6
port 11 n
rlabel metal3 161061 16808 161861 16928 1 Bit5
port 12 n
rlabel metal3 161061 18576 161861 18696 1 Bit4
port 13 n
rlabel metal3 161061 20344 161861 20464 1 Bit3
port 14 n
rlabel metal3 161061 22112 161861 22232 1 Bit2
port 15 n
rlabel metal3 161061 23880 161861 24000 1 Bit1
port 16 n
rlabel metal3 161061 29184 161861 29304 1 RESET
port 17 n
<< end >>
