magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -386 144812 386 144840
rect -386 140578 302 144812
rect 366 140578 386 144812
rect -386 140550 386 140578
rect -386 140282 386 140310
rect -386 136048 302 140282
rect 366 136048 386 140282
rect -386 136020 386 136048
rect -386 135752 386 135780
rect -386 131518 302 135752
rect 366 131518 386 135752
rect -386 131490 386 131518
rect -386 131222 386 131250
rect -386 126988 302 131222
rect 366 126988 386 131222
rect -386 126960 386 126988
rect -386 126692 386 126720
rect -386 122458 302 126692
rect 366 122458 386 126692
rect -386 122430 386 122458
rect -386 122162 386 122190
rect -386 117928 302 122162
rect 366 117928 386 122162
rect -386 117900 386 117928
rect -386 117632 386 117660
rect -386 113398 302 117632
rect 366 113398 386 117632
rect -386 113370 386 113398
rect -386 113102 386 113130
rect -386 108868 302 113102
rect 366 108868 386 113102
rect -386 108840 386 108868
rect -386 108572 386 108600
rect -386 104338 302 108572
rect 366 104338 386 108572
rect -386 104310 386 104338
rect -386 104042 386 104070
rect -386 99808 302 104042
rect 366 99808 386 104042
rect -386 99780 386 99808
rect -386 99512 386 99540
rect -386 95278 302 99512
rect 366 95278 386 99512
rect -386 95250 386 95278
rect -386 94982 386 95010
rect -386 90748 302 94982
rect 366 90748 386 94982
rect -386 90720 386 90748
rect -386 90452 386 90480
rect -386 86218 302 90452
rect 366 86218 386 90452
rect -386 86190 386 86218
rect -386 85922 386 85950
rect -386 81688 302 85922
rect 366 81688 386 85922
rect -386 81660 386 81688
rect -386 81392 386 81420
rect -386 77158 302 81392
rect 366 77158 386 81392
rect -386 77130 386 77158
rect -386 76862 386 76890
rect -386 72628 302 76862
rect 366 72628 386 76862
rect -386 72600 386 72628
rect -386 72332 386 72360
rect -386 68098 302 72332
rect 366 68098 386 72332
rect -386 68070 386 68098
rect -386 67802 386 67830
rect -386 63568 302 67802
rect 366 63568 386 67802
rect -386 63540 386 63568
rect -386 63272 386 63300
rect -386 59038 302 63272
rect 366 59038 386 63272
rect -386 59010 386 59038
rect -386 58742 386 58770
rect -386 54508 302 58742
rect 366 54508 386 58742
rect -386 54480 386 54508
rect -386 54212 386 54240
rect -386 49978 302 54212
rect 366 49978 386 54212
rect -386 49950 386 49978
rect -386 49682 386 49710
rect -386 45448 302 49682
rect 366 45448 386 49682
rect -386 45420 386 45448
rect -386 45152 386 45180
rect -386 40918 302 45152
rect 366 40918 386 45152
rect -386 40890 386 40918
rect -386 40622 386 40650
rect -386 36388 302 40622
rect 366 36388 386 40622
rect -386 36360 386 36388
rect -386 36092 386 36120
rect -386 31858 302 36092
rect 366 31858 386 36092
rect -386 31830 386 31858
rect -386 31562 386 31590
rect -386 27328 302 31562
rect 366 27328 386 31562
rect -386 27300 386 27328
rect -386 27032 386 27060
rect -386 22798 302 27032
rect 366 22798 386 27032
rect -386 22770 386 22798
rect -386 22502 386 22530
rect -386 18268 302 22502
rect 366 18268 386 22502
rect -386 18240 386 18268
rect -386 17972 386 18000
rect -386 13738 302 17972
rect 366 13738 386 17972
rect -386 13710 386 13738
rect -386 13442 386 13470
rect -386 9208 302 13442
rect 366 9208 386 13442
rect -386 9180 386 9208
rect -386 8912 386 8940
rect -386 4678 302 8912
rect 366 4678 386 8912
rect -386 4650 386 4678
rect -386 4382 386 4410
rect -386 148 302 4382
rect 366 148 386 4382
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -4382 302 -148
rect 366 -4382 386 -148
rect -386 -4410 386 -4382
rect -386 -4678 386 -4650
rect -386 -8912 302 -4678
rect 366 -8912 386 -4678
rect -386 -8940 386 -8912
rect -386 -9208 386 -9180
rect -386 -13442 302 -9208
rect 366 -13442 386 -9208
rect -386 -13470 386 -13442
rect -386 -13738 386 -13710
rect -386 -17972 302 -13738
rect 366 -17972 386 -13738
rect -386 -18000 386 -17972
rect -386 -18268 386 -18240
rect -386 -22502 302 -18268
rect 366 -22502 386 -18268
rect -386 -22530 386 -22502
rect -386 -22798 386 -22770
rect -386 -27032 302 -22798
rect 366 -27032 386 -22798
rect -386 -27060 386 -27032
rect -386 -27328 386 -27300
rect -386 -31562 302 -27328
rect 366 -31562 386 -27328
rect -386 -31590 386 -31562
rect -386 -31858 386 -31830
rect -386 -36092 302 -31858
rect 366 -36092 386 -31858
rect -386 -36120 386 -36092
rect -386 -36388 386 -36360
rect -386 -40622 302 -36388
rect 366 -40622 386 -36388
rect -386 -40650 386 -40622
rect -386 -40918 386 -40890
rect -386 -45152 302 -40918
rect 366 -45152 386 -40918
rect -386 -45180 386 -45152
rect -386 -45448 386 -45420
rect -386 -49682 302 -45448
rect 366 -49682 386 -45448
rect -386 -49710 386 -49682
rect -386 -49978 386 -49950
rect -386 -54212 302 -49978
rect 366 -54212 386 -49978
rect -386 -54240 386 -54212
rect -386 -54508 386 -54480
rect -386 -58742 302 -54508
rect 366 -58742 386 -54508
rect -386 -58770 386 -58742
rect -386 -59038 386 -59010
rect -386 -63272 302 -59038
rect 366 -63272 386 -59038
rect -386 -63300 386 -63272
rect -386 -63568 386 -63540
rect -386 -67802 302 -63568
rect 366 -67802 386 -63568
rect -386 -67830 386 -67802
rect -386 -68098 386 -68070
rect -386 -72332 302 -68098
rect 366 -72332 386 -68098
rect -386 -72360 386 -72332
rect -386 -72628 386 -72600
rect -386 -76862 302 -72628
rect 366 -76862 386 -72628
rect -386 -76890 386 -76862
rect -386 -77158 386 -77130
rect -386 -81392 302 -77158
rect 366 -81392 386 -77158
rect -386 -81420 386 -81392
rect -386 -81688 386 -81660
rect -386 -85922 302 -81688
rect 366 -85922 386 -81688
rect -386 -85950 386 -85922
rect -386 -86218 386 -86190
rect -386 -90452 302 -86218
rect 366 -90452 386 -86218
rect -386 -90480 386 -90452
rect -386 -90748 386 -90720
rect -386 -94982 302 -90748
rect 366 -94982 386 -90748
rect -386 -95010 386 -94982
rect -386 -95278 386 -95250
rect -386 -99512 302 -95278
rect 366 -99512 386 -95278
rect -386 -99540 386 -99512
rect -386 -99808 386 -99780
rect -386 -104042 302 -99808
rect 366 -104042 386 -99808
rect -386 -104070 386 -104042
rect -386 -104338 386 -104310
rect -386 -108572 302 -104338
rect 366 -108572 386 -104338
rect -386 -108600 386 -108572
rect -386 -108868 386 -108840
rect -386 -113102 302 -108868
rect 366 -113102 386 -108868
rect -386 -113130 386 -113102
rect -386 -113398 386 -113370
rect -386 -117632 302 -113398
rect 366 -117632 386 -113398
rect -386 -117660 386 -117632
rect -386 -117928 386 -117900
rect -386 -122162 302 -117928
rect 366 -122162 386 -117928
rect -386 -122190 386 -122162
rect -386 -122458 386 -122430
rect -386 -126692 302 -122458
rect 366 -126692 386 -122458
rect -386 -126720 386 -126692
rect -386 -126988 386 -126960
rect -386 -131222 302 -126988
rect 366 -131222 386 -126988
rect -386 -131250 386 -131222
rect -386 -131518 386 -131490
rect -386 -135752 302 -131518
rect 366 -135752 386 -131518
rect -386 -135780 386 -135752
rect -386 -136048 386 -136020
rect -386 -140282 302 -136048
rect 366 -140282 386 -136048
rect -386 -140310 386 -140282
rect -386 -140578 386 -140550
rect -386 -144812 302 -140578
rect 366 -144812 386 -140578
rect -386 -144840 386 -144812
<< via3 >>
rect 302 140578 366 144812
rect 302 136048 366 140282
rect 302 131518 366 135752
rect 302 126988 366 131222
rect 302 122458 366 126692
rect 302 117928 366 122162
rect 302 113398 366 117632
rect 302 108868 366 113102
rect 302 104338 366 108572
rect 302 99808 366 104042
rect 302 95278 366 99512
rect 302 90748 366 94982
rect 302 86218 366 90452
rect 302 81688 366 85922
rect 302 77158 366 81392
rect 302 72628 366 76862
rect 302 68098 366 72332
rect 302 63568 366 67802
rect 302 59038 366 63272
rect 302 54508 366 58742
rect 302 49978 366 54212
rect 302 45448 366 49682
rect 302 40918 366 45152
rect 302 36388 366 40622
rect 302 31858 366 36092
rect 302 27328 366 31562
rect 302 22798 366 27032
rect 302 18268 366 22502
rect 302 13738 366 17972
rect 302 9208 366 13442
rect 302 4678 366 8912
rect 302 148 366 4382
rect 302 -4382 366 -148
rect 302 -8912 366 -4678
rect 302 -13442 366 -9208
rect 302 -17972 366 -13738
rect 302 -22502 366 -18268
rect 302 -27032 366 -22798
rect 302 -31562 366 -27328
rect 302 -36092 366 -31858
rect 302 -40622 366 -36388
rect 302 -45152 366 -40918
rect 302 -49682 366 -45448
rect 302 -54212 366 -49978
rect 302 -58742 366 -54508
rect 302 -63272 366 -59038
rect 302 -67802 366 -63568
rect 302 -72332 366 -68098
rect 302 -76862 366 -72628
rect 302 -81392 366 -77158
rect 302 -85922 366 -81688
rect 302 -90452 366 -86218
rect 302 -94982 366 -90748
rect 302 -99512 366 -95278
rect 302 -104042 366 -99808
rect 302 -108572 366 -104338
rect 302 -113102 366 -108868
rect 302 -117632 366 -113398
rect 302 -122162 366 -117928
rect 302 -126692 366 -122458
rect 302 -131222 366 -126988
rect 302 -135752 366 -131518
rect 302 -140282 366 -136048
rect 302 -144812 366 -140578
<< mimcap >>
rect -346 144760 54 144800
rect -346 140630 -306 144760
rect 14 140630 54 144760
rect -346 140590 54 140630
rect -346 140230 54 140270
rect -346 136100 -306 140230
rect 14 136100 54 140230
rect -346 136060 54 136100
rect -346 135700 54 135740
rect -346 131570 -306 135700
rect 14 131570 54 135700
rect -346 131530 54 131570
rect -346 131170 54 131210
rect -346 127040 -306 131170
rect 14 127040 54 131170
rect -346 127000 54 127040
rect -346 126640 54 126680
rect -346 122510 -306 126640
rect 14 122510 54 126640
rect -346 122470 54 122510
rect -346 122110 54 122150
rect -346 117980 -306 122110
rect 14 117980 54 122110
rect -346 117940 54 117980
rect -346 117580 54 117620
rect -346 113450 -306 117580
rect 14 113450 54 117580
rect -346 113410 54 113450
rect -346 113050 54 113090
rect -346 108920 -306 113050
rect 14 108920 54 113050
rect -346 108880 54 108920
rect -346 108520 54 108560
rect -346 104390 -306 108520
rect 14 104390 54 108520
rect -346 104350 54 104390
rect -346 103990 54 104030
rect -346 99860 -306 103990
rect 14 99860 54 103990
rect -346 99820 54 99860
rect -346 99460 54 99500
rect -346 95330 -306 99460
rect 14 95330 54 99460
rect -346 95290 54 95330
rect -346 94930 54 94970
rect -346 90800 -306 94930
rect 14 90800 54 94930
rect -346 90760 54 90800
rect -346 90400 54 90440
rect -346 86270 -306 90400
rect 14 86270 54 90400
rect -346 86230 54 86270
rect -346 85870 54 85910
rect -346 81740 -306 85870
rect 14 81740 54 85870
rect -346 81700 54 81740
rect -346 81340 54 81380
rect -346 77210 -306 81340
rect 14 77210 54 81340
rect -346 77170 54 77210
rect -346 76810 54 76850
rect -346 72680 -306 76810
rect 14 72680 54 76810
rect -346 72640 54 72680
rect -346 72280 54 72320
rect -346 68150 -306 72280
rect 14 68150 54 72280
rect -346 68110 54 68150
rect -346 67750 54 67790
rect -346 63620 -306 67750
rect 14 63620 54 67750
rect -346 63580 54 63620
rect -346 63220 54 63260
rect -346 59090 -306 63220
rect 14 59090 54 63220
rect -346 59050 54 59090
rect -346 58690 54 58730
rect -346 54560 -306 58690
rect 14 54560 54 58690
rect -346 54520 54 54560
rect -346 54160 54 54200
rect -346 50030 -306 54160
rect 14 50030 54 54160
rect -346 49990 54 50030
rect -346 49630 54 49670
rect -346 45500 -306 49630
rect 14 45500 54 49630
rect -346 45460 54 45500
rect -346 45100 54 45140
rect -346 40970 -306 45100
rect 14 40970 54 45100
rect -346 40930 54 40970
rect -346 40570 54 40610
rect -346 36440 -306 40570
rect 14 36440 54 40570
rect -346 36400 54 36440
rect -346 36040 54 36080
rect -346 31910 -306 36040
rect 14 31910 54 36040
rect -346 31870 54 31910
rect -346 31510 54 31550
rect -346 27380 -306 31510
rect 14 27380 54 31510
rect -346 27340 54 27380
rect -346 26980 54 27020
rect -346 22850 -306 26980
rect 14 22850 54 26980
rect -346 22810 54 22850
rect -346 22450 54 22490
rect -346 18320 -306 22450
rect 14 18320 54 22450
rect -346 18280 54 18320
rect -346 17920 54 17960
rect -346 13790 -306 17920
rect 14 13790 54 17920
rect -346 13750 54 13790
rect -346 13390 54 13430
rect -346 9260 -306 13390
rect 14 9260 54 13390
rect -346 9220 54 9260
rect -346 8860 54 8900
rect -346 4730 -306 8860
rect 14 4730 54 8860
rect -346 4690 54 4730
rect -346 4330 54 4370
rect -346 200 -306 4330
rect 14 200 54 4330
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -4330 -306 -200
rect 14 -4330 54 -200
rect -346 -4370 54 -4330
rect -346 -4730 54 -4690
rect -346 -8860 -306 -4730
rect 14 -8860 54 -4730
rect -346 -8900 54 -8860
rect -346 -9260 54 -9220
rect -346 -13390 -306 -9260
rect 14 -13390 54 -9260
rect -346 -13430 54 -13390
rect -346 -13790 54 -13750
rect -346 -17920 -306 -13790
rect 14 -17920 54 -13790
rect -346 -17960 54 -17920
rect -346 -18320 54 -18280
rect -346 -22450 -306 -18320
rect 14 -22450 54 -18320
rect -346 -22490 54 -22450
rect -346 -22850 54 -22810
rect -346 -26980 -306 -22850
rect 14 -26980 54 -22850
rect -346 -27020 54 -26980
rect -346 -27380 54 -27340
rect -346 -31510 -306 -27380
rect 14 -31510 54 -27380
rect -346 -31550 54 -31510
rect -346 -31910 54 -31870
rect -346 -36040 -306 -31910
rect 14 -36040 54 -31910
rect -346 -36080 54 -36040
rect -346 -36440 54 -36400
rect -346 -40570 -306 -36440
rect 14 -40570 54 -36440
rect -346 -40610 54 -40570
rect -346 -40970 54 -40930
rect -346 -45100 -306 -40970
rect 14 -45100 54 -40970
rect -346 -45140 54 -45100
rect -346 -45500 54 -45460
rect -346 -49630 -306 -45500
rect 14 -49630 54 -45500
rect -346 -49670 54 -49630
rect -346 -50030 54 -49990
rect -346 -54160 -306 -50030
rect 14 -54160 54 -50030
rect -346 -54200 54 -54160
rect -346 -54560 54 -54520
rect -346 -58690 -306 -54560
rect 14 -58690 54 -54560
rect -346 -58730 54 -58690
rect -346 -59090 54 -59050
rect -346 -63220 -306 -59090
rect 14 -63220 54 -59090
rect -346 -63260 54 -63220
rect -346 -63620 54 -63580
rect -346 -67750 -306 -63620
rect 14 -67750 54 -63620
rect -346 -67790 54 -67750
rect -346 -68150 54 -68110
rect -346 -72280 -306 -68150
rect 14 -72280 54 -68150
rect -346 -72320 54 -72280
rect -346 -72680 54 -72640
rect -346 -76810 -306 -72680
rect 14 -76810 54 -72680
rect -346 -76850 54 -76810
rect -346 -77210 54 -77170
rect -346 -81340 -306 -77210
rect 14 -81340 54 -77210
rect -346 -81380 54 -81340
rect -346 -81740 54 -81700
rect -346 -85870 -306 -81740
rect 14 -85870 54 -81740
rect -346 -85910 54 -85870
rect -346 -86270 54 -86230
rect -346 -90400 -306 -86270
rect 14 -90400 54 -86270
rect -346 -90440 54 -90400
rect -346 -90800 54 -90760
rect -346 -94930 -306 -90800
rect 14 -94930 54 -90800
rect -346 -94970 54 -94930
rect -346 -95330 54 -95290
rect -346 -99460 -306 -95330
rect 14 -99460 54 -95330
rect -346 -99500 54 -99460
rect -346 -99860 54 -99820
rect -346 -103990 -306 -99860
rect 14 -103990 54 -99860
rect -346 -104030 54 -103990
rect -346 -104390 54 -104350
rect -346 -108520 -306 -104390
rect 14 -108520 54 -104390
rect -346 -108560 54 -108520
rect -346 -108920 54 -108880
rect -346 -113050 -306 -108920
rect 14 -113050 54 -108920
rect -346 -113090 54 -113050
rect -346 -113450 54 -113410
rect -346 -117580 -306 -113450
rect 14 -117580 54 -113450
rect -346 -117620 54 -117580
rect -346 -117980 54 -117940
rect -346 -122110 -306 -117980
rect 14 -122110 54 -117980
rect -346 -122150 54 -122110
rect -346 -122510 54 -122470
rect -346 -126640 -306 -122510
rect 14 -126640 54 -122510
rect -346 -126680 54 -126640
rect -346 -127040 54 -127000
rect -346 -131170 -306 -127040
rect 14 -131170 54 -127040
rect -346 -131210 54 -131170
rect -346 -131570 54 -131530
rect -346 -135700 -306 -131570
rect 14 -135700 54 -131570
rect -346 -135740 54 -135700
rect -346 -136100 54 -136060
rect -346 -140230 -306 -136100
rect 14 -140230 54 -136100
rect -346 -140270 54 -140230
rect -346 -140630 54 -140590
rect -346 -144760 -306 -140630
rect 14 -144760 54 -140630
rect -346 -144800 54 -144760
<< mimcapcontact >>
rect -306 140630 14 144760
rect -306 136100 14 140230
rect -306 131570 14 135700
rect -306 127040 14 131170
rect -306 122510 14 126640
rect -306 117980 14 122110
rect -306 113450 14 117580
rect -306 108920 14 113050
rect -306 104390 14 108520
rect -306 99860 14 103990
rect -306 95330 14 99460
rect -306 90800 14 94930
rect -306 86270 14 90400
rect -306 81740 14 85870
rect -306 77210 14 81340
rect -306 72680 14 76810
rect -306 68150 14 72280
rect -306 63620 14 67750
rect -306 59090 14 63220
rect -306 54560 14 58690
rect -306 50030 14 54160
rect -306 45500 14 49630
rect -306 40970 14 45100
rect -306 36440 14 40570
rect -306 31910 14 36040
rect -306 27380 14 31510
rect -306 22850 14 26980
rect -306 18320 14 22450
rect -306 13790 14 17920
rect -306 9260 14 13390
rect -306 4730 14 8860
rect -306 200 14 4330
rect -306 -4330 14 -200
rect -306 -8860 14 -4730
rect -306 -13390 14 -9260
rect -306 -17920 14 -13790
rect -306 -22450 14 -18320
rect -306 -26980 14 -22850
rect -306 -31510 14 -27380
rect -306 -36040 14 -31910
rect -306 -40570 14 -36440
rect -306 -45100 14 -40970
rect -306 -49630 14 -45500
rect -306 -54160 14 -50030
rect -306 -58690 14 -54560
rect -306 -63220 14 -59090
rect -306 -67750 14 -63620
rect -306 -72280 14 -68150
rect -306 -76810 14 -72680
rect -306 -81340 14 -77210
rect -306 -85870 14 -81740
rect -306 -90400 14 -86270
rect -306 -94930 14 -90800
rect -306 -99460 14 -95330
rect -306 -103990 14 -99860
rect -306 -108520 14 -104390
rect -306 -113050 14 -108920
rect -306 -117580 14 -113450
rect -306 -122110 14 -117980
rect -306 -126640 14 -122510
rect -306 -131170 14 -127040
rect -306 -135700 14 -131570
rect -306 -140230 14 -136100
rect -306 -144760 14 -140630
<< metal4 >>
rect -198 144761 -94 144960
rect 282 144812 386 144960
rect -307 144760 15 144761
rect -307 140630 -306 144760
rect 14 140630 15 144760
rect -307 140629 15 140630
rect -198 140231 -94 140629
rect 282 140578 302 144812
rect 366 140578 386 144812
rect 282 140282 386 140578
rect -307 140230 15 140231
rect -307 136100 -306 140230
rect 14 136100 15 140230
rect -307 136099 15 136100
rect -198 135701 -94 136099
rect 282 136048 302 140282
rect 366 136048 386 140282
rect 282 135752 386 136048
rect -307 135700 15 135701
rect -307 131570 -306 135700
rect 14 131570 15 135700
rect -307 131569 15 131570
rect -198 131171 -94 131569
rect 282 131518 302 135752
rect 366 131518 386 135752
rect 282 131222 386 131518
rect -307 131170 15 131171
rect -307 127040 -306 131170
rect 14 127040 15 131170
rect -307 127039 15 127040
rect -198 126641 -94 127039
rect 282 126988 302 131222
rect 366 126988 386 131222
rect 282 126692 386 126988
rect -307 126640 15 126641
rect -307 122510 -306 126640
rect 14 122510 15 126640
rect -307 122509 15 122510
rect -198 122111 -94 122509
rect 282 122458 302 126692
rect 366 122458 386 126692
rect 282 122162 386 122458
rect -307 122110 15 122111
rect -307 117980 -306 122110
rect 14 117980 15 122110
rect -307 117979 15 117980
rect -198 117581 -94 117979
rect 282 117928 302 122162
rect 366 117928 386 122162
rect 282 117632 386 117928
rect -307 117580 15 117581
rect -307 113450 -306 117580
rect 14 113450 15 117580
rect -307 113449 15 113450
rect -198 113051 -94 113449
rect 282 113398 302 117632
rect 366 113398 386 117632
rect 282 113102 386 113398
rect -307 113050 15 113051
rect -307 108920 -306 113050
rect 14 108920 15 113050
rect -307 108919 15 108920
rect -198 108521 -94 108919
rect 282 108868 302 113102
rect 366 108868 386 113102
rect 282 108572 386 108868
rect -307 108520 15 108521
rect -307 104390 -306 108520
rect 14 104390 15 108520
rect -307 104389 15 104390
rect -198 103991 -94 104389
rect 282 104338 302 108572
rect 366 104338 386 108572
rect 282 104042 386 104338
rect -307 103990 15 103991
rect -307 99860 -306 103990
rect 14 99860 15 103990
rect -307 99859 15 99860
rect -198 99461 -94 99859
rect 282 99808 302 104042
rect 366 99808 386 104042
rect 282 99512 386 99808
rect -307 99460 15 99461
rect -307 95330 -306 99460
rect 14 95330 15 99460
rect -307 95329 15 95330
rect -198 94931 -94 95329
rect 282 95278 302 99512
rect 366 95278 386 99512
rect 282 94982 386 95278
rect -307 94930 15 94931
rect -307 90800 -306 94930
rect 14 90800 15 94930
rect -307 90799 15 90800
rect -198 90401 -94 90799
rect 282 90748 302 94982
rect 366 90748 386 94982
rect 282 90452 386 90748
rect -307 90400 15 90401
rect -307 86270 -306 90400
rect 14 86270 15 90400
rect -307 86269 15 86270
rect -198 85871 -94 86269
rect 282 86218 302 90452
rect 366 86218 386 90452
rect 282 85922 386 86218
rect -307 85870 15 85871
rect -307 81740 -306 85870
rect 14 81740 15 85870
rect -307 81739 15 81740
rect -198 81341 -94 81739
rect 282 81688 302 85922
rect 366 81688 386 85922
rect 282 81392 386 81688
rect -307 81340 15 81341
rect -307 77210 -306 81340
rect 14 77210 15 81340
rect -307 77209 15 77210
rect -198 76811 -94 77209
rect 282 77158 302 81392
rect 366 77158 386 81392
rect 282 76862 386 77158
rect -307 76810 15 76811
rect -307 72680 -306 76810
rect 14 72680 15 76810
rect -307 72679 15 72680
rect -198 72281 -94 72679
rect 282 72628 302 76862
rect 366 72628 386 76862
rect 282 72332 386 72628
rect -307 72280 15 72281
rect -307 68150 -306 72280
rect 14 68150 15 72280
rect -307 68149 15 68150
rect -198 67751 -94 68149
rect 282 68098 302 72332
rect 366 68098 386 72332
rect 282 67802 386 68098
rect -307 67750 15 67751
rect -307 63620 -306 67750
rect 14 63620 15 67750
rect -307 63619 15 63620
rect -198 63221 -94 63619
rect 282 63568 302 67802
rect 366 63568 386 67802
rect 282 63272 386 63568
rect -307 63220 15 63221
rect -307 59090 -306 63220
rect 14 59090 15 63220
rect -307 59089 15 59090
rect -198 58691 -94 59089
rect 282 59038 302 63272
rect 366 59038 386 63272
rect 282 58742 386 59038
rect -307 58690 15 58691
rect -307 54560 -306 58690
rect 14 54560 15 58690
rect -307 54559 15 54560
rect -198 54161 -94 54559
rect 282 54508 302 58742
rect 366 54508 386 58742
rect 282 54212 386 54508
rect -307 54160 15 54161
rect -307 50030 -306 54160
rect 14 50030 15 54160
rect -307 50029 15 50030
rect -198 49631 -94 50029
rect 282 49978 302 54212
rect 366 49978 386 54212
rect 282 49682 386 49978
rect -307 49630 15 49631
rect -307 45500 -306 49630
rect 14 45500 15 49630
rect -307 45499 15 45500
rect -198 45101 -94 45499
rect 282 45448 302 49682
rect 366 45448 386 49682
rect 282 45152 386 45448
rect -307 45100 15 45101
rect -307 40970 -306 45100
rect 14 40970 15 45100
rect -307 40969 15 40970
rect -198 40571 -94 40969
rect 282 40918 302 45152
rect 366 40918 386 45152
rect 282 40622 386 40918
rect -307 40570 15 40571
rect -307 36440 -306 40570
rect 14 36440 15 40570
rect -307 36439 15 36440
rect -198 36041 -94 36439
rect 282 36388 302 40622
rect 366 36388 386 40622
rect 282 36092 386 36388
rect -307 36040 15 36041
rect -307 31910 -306 36040
rect 14 31910 15 36040
rect -307 31909 15 31910
rect -198 31511 -94 31909
rect 282 31858 302 36092
rect 366 31858 386 36092
rect 282 31562 386 31858
rect -307 31510 15 31511
rect -307 27380 -306 31510
rect 14 27380 15 31510
rect -307 27379 15 27380
rect -198 26981 -94 27379
rect 282 27328 302 31562
rect 366 27328 386 31562
rect 282 27032 386 27328
rect -307 26980 15 26981
rect -307 22850 -306 26980
rect 14 22850 15 26980
rect -307 22849 15 22850
rect -198 22451 -94 22849
rect 282 22798 302 27032
rect 366 22798 386 27032
rect 282 22502 386 22798
rect -307 22450 15 22451
rect -307 18320 -306 22450
rect 14 18320 15 22450
rect -307 18319 15 18320
rect -198 17921 -94 18319
rect 282 18268 302 22502
rect 366 18268 386 22502
rect 282 17972 386 18268
rect -307 17920 15 17921
rect -307 13790 -306 17920
rect 14 13790 15 17920
rect -307 13789 15 13790
rect -198 13391 -94 13789
rect 282 13738 302 17972
rect 366 13738 386 17972
rect 282 13442 386 13738
rect -307 13390 15 13391
rect -307 9260 -306 13390
rect 14 9260 15 13390
rect -307 9259 15 9260
rect -198 8861 -94 9259
rect 282 9208 302 13442
rect 366 9208 386 13442
rect 282 8912 386 9208
rect -307 8860 15 8861
rect -307 4730 -306 8860
rect 14 4730 15 8860
rect -307 4729 15 4730
rect -198 4331 -94 4729
rect 282 4678 302 8912
rect 366 4678 386 8912
rect 282 4382 386 4678
rect -307 4330 15 4331
rect -307 200 -306 4330
rect 14 200 15 4330
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 4382
rect 366 148 386 4382
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -4330 -306 -200
rect 14 -4330 15 -200
rect -307 -4331 15 -4330
rect -198 -4729 -94 -4331
rect 282 -4382 302 -148
rect 366 -4382 386 -148
rect 282 -4678 386 -4382
rect -307 -4730 15 -4729
rect -307 -8860 -306 -4730
rect 14 -8860 15 -4730
rect -307 -8861 15 -8860
rect -198 -9259 -94 -8861
rect 282 -8912 302 -4678
rect 366 -8912 386 -4678
rect 282 -9208 386 -8912
rect -307 -9260 15 -9259
rect -307 -13390 -306 -9260
rect 14 -13390 15 -9260
rect -307 -13391 15 -13390
rect -198 -13789 -94 -13391
rect 282 -13442 302 -9208
rect 366 -13442 386 -9208
rect 282 -13738 386 -13442
rect -307 -13790 15 -13789
rect -307 -17920 -306 -13790
rect 14 -17920 15 -13790
rect -307 -17921 15 -17920
rect -198 -18319 -94 -17921
rect 282 -17972 302 -13738
rect 366 -17972 386 -13738
rect 282 -18268 386 -17972
rect -307 -18320 15 -18319
rect -307 -22450 -306 -18320
rect 14 -22450 15 -18320
rect -307 -22451 15 -22450
rect -198 -22849 -94 -22451
rect 282 -22502 302 -18268
rect 366 -22502 386 -18268
rect 282 -22798 386 -22502
rect -307 -22850 15 -22849
rect -307 -26980 -306 -22850
rect 14 -26980 15 -22850
rect -307 -26981 15 -26980
rect -198 -27379 -94 -26981
rect 282 -27032 302 -22798
rect 366 -27032 386 -22798
rect 282 -27328 386 -27032
rect -307 -27380 15 -27379
rect -307 -31510 -306 -27380
rect 14 -31510 15 -27380
rect -307 -31511 15 -31510
rect -198 -31909 -94 -31511
rect 282 -31562 302 -27328
rect 366 -31562 386 -27328
rect 282 -31858 386 -31562
rect -307 -31910 15 -31909
rect -307 -36040 -306 -31910
rect 14 -36040 15 -31910
rect -307 -36041 15 -36040
rect -198 -36439 -94 -36041
rect 282 -36092 302 -31858
rect 366 -36092 386 -31858
rect 282 -36388 386 -36092
rect -307 -36440 15 -36439
rect -307 -40570 -306 -36440
rect 14 -40570 15 -36440
rect -307 -40571 15 -40570
rect -198 -40969 -94 -40571
rect 282 -40622 302 -36388
rect 366 -40622 386 -36388
rect 282 -40918 386 -40622
rect -307 -40970 15 -40969
rect -307 -45100 -306 -40970
rect 14 -45100 15 -40970
rect -307 -45101 15 -45100
rect -198 -45499 -94 -45101
rect 282 -45152 302 -40918
rect 366 -45152 386 -40918
rect 282 -45448 386 -45152
rect -307 -45500 15 -45499
rect -307 -49630 -306 -45500
rect 14 -49630 15 -45500
rect -307 -49631 15 -49630
rect -198 -50029 -94 -49631
rect 282 -49682 302 -45448
rect 366 -49682 386 -45448
rect 282 -49978 386 -49682
rect -307 -50030 15 -50029
rect -307 -54160 -306 -50030
rect 14 -54160 15 -50030
rect -307 -54161 15 -54160
rect -198 -54559 -94 -54161
rect 282 -54212 302 -49978
rect 366 -54212 386 -49978
rect 282 -54508 386 -54212
rect -307 -54560 15 -54559
rect -307 -58690 -306 -54560
rect 14 -58690 15 -54560
rect -307 -58691 15 -58690
rect -198 -59089 -94 -58691
rect 282 -58742 302 -54508
rect 366 -58742 386 -54508
rect 282 -59038 386 -58742
rect -307 -59090 15 -59089
rect -307 -63220 -306 -59090
rect 14 -63220 15 -59090
rect -307 -63221 15 -63220
rect -198 -63619 -94 -63221
rect 282 -63272 302 -59038
rect 366 -63272 386 -59038
rect 282 -63568 386 -63272
rect -307 -63620 15 -63619
rect -307 -67750 -306 -63620
rect 14 -67750 15 -63620
rect -307 -67751 15 -67750
rect -198 -68149 -94 -67751
rect 282 -67802 302 -63568
rect 366 -67802 386 -63568
rect 282 -68098 386 -67802
rect -307 -68150 15 -68149
rect -307 -72280 -306 -68150
rect 14 -72280 15 -68150
rect -307 -72281 15 -72280
rect -198 -72679 -94 -72281
rect 282 -72332 302 -68098
rect 366 -72332 386 -68098
rect 282 -72628 386 -72332
rect -307 -72680 15 -72679
rect -307 -76810 -306 -72680
rect 14 -76810 15 -72680
rect -307 -76811 15 -76810
rect -198 -77209 -94 -76811
rect 282 -76862 302 -72628
rect 366 -76862 386 -72628
rect 282 -77158 386 -76862
rect -307 -77210 15 -77209
rect -307 -81340 -306 -77210
rect 14 -81340 15 -77210
rect -307 -81341 15 -81340
rect -198 -81739 -94 -81341
rect 282 -81392 302 -77158
rect 366 -81392 386 -77158
rect 282 -81688 386 -81392
rect -307 -81740 15 -81739
rect -307 -85870 -306 -81740
rect 14 -85870 15 -81740
rect -307 -85871 15 -85870
rect -198 -86269 -94 -85871
rect 282 -85922 302 -81688
rect 366 -85922 386 -81688
rect 282 -86218 386 -85922
rect -307 -86270 15 -86269
rect -307 -90400 -306 -86270
rect 14 -90400 15 -86270
rect -307 -90401 15 -90400
rect -198 -90799 -94 -90401
rect 282 -90452 302 -86218
rect 366 -90452 386 -86218
rect 282 -90748 386 -90452
rect -307 -90800 15 -90799
rect -307 -94930 -306 -90800
rect 14 -94930 15 -90800
rect -307 -94931 15 -94930
rect -198 -95329 -94 -94931
rect 282 -94982 302 -90748
rect 366 -94982 386 -90748
rect 282 -95278 386 -94982
rect -307 -95330 15 -95329
rect -307 -99460 -306 -95330
rect 14 -99460 15 -95330
rect -307 -99461 15 -99460
rect -198 -99859 -94 -99461
rect 282 -99512 302 -95278
rect 366 -99512 386 -95278
rect 282 -99808 386 -99512
rect -307 -99860 15 -99859
rect -307 -103990 -306 -99860
rect 14 -103990 15 -99860
rect -307 -103991 15 -103990
rect -198 -104389 -94 -103991
rect 282 -104042 302 -99808
rect 366 -104042 386 -99808
rect 282 -104338 386 -104042
rect -307 -104390 15 -104389
rect -307 -108520 -306 -104390
rect 14 -108520 15 -104390
rect -307 -108521 15 -108520
rect -198 -108919 -94 -108521
rect 282 -108572 302 -104338
rect 366 -108572 386 -104338
rect 282 -108868 386 -108572
rect -307 -108920 15 -108919
rect -307 -113050 -306 -108920
rect 14 -113050 15 -108920
rect -307 -113051 15 -113050
rect -198 -113449 -94 -113051
rect 282 -113102 302 -108868
rect 366 -113102 386 -108868
rect 282 -113398 386 -113102
rect -307 -113450 15 -113449
rect -307 -117580 -306 -113450
rect 14 -117580 15 -113450
rect -307 -117581 15 -117580
rect -198 -117979 -94 -117581
rect 282 -117632 302 -113398
rect 366 -117632 386 -113398
rect 282 -117928 386 -117632
rect -307 -117980 15 -117979
rect -307 -122110 -306 -117980
rect 14 -122110 15 -117980
rect -307 -122111 15 -122110
rect -198 -122509 -94 -122111
rect 282 -122162 302 -117928
rect 366 -122162 386 -117928
rect 282 -122458 386 -122162
rect -307 -122510 15 -122509
rect -307 -126640 -306 -122510
rect 14 -126640 15 -122510
rect -307 -126641 15 -126640
rect -198 -127039 -94 -126641
rect 282 -126692 302 -122458
rect 366 -126692 386 -122458
rect 282 -126988 386 -126692
rect -307 -127040 15 -127039
rect -307 -131170 -306 -127040
rect 14 -131170 15 -127040
rect -307 -131171 15 -131170
rect -198 -131569 -94 -131171
rect 282 -131222 302 -126988
rect 366 -131222 386 -126988
rect 282 -131518 386 -131222
rect -307 -131570 15 -131569
rect -307 -135700 -306 -131570
rect 14 -135700 15 -131570
rect -307 -135701 15 -135700
rect -198 -136099 -94 -135701
rect 282 -135752 302 -131518
rect 366 -135752 386 -131518
rect 282 -136048 386 -135752
rect -307 -136100 15 -136099
rect -307 -140230 -306 -136100
rect 14 -140230 15 -136100
rect -307 -140231 15 -140230
rect -198 -140629 -94 -140231
rect 282 -140282 302 -136048
rect 366 -140282 386 -136048
rect 282 -140578 386 -140282
rect -307 -140630 15 -140629
rect -307 -144760 -306 -140630
rect 14 -144760 15 -140630
rect -307 -144761 15 -144760
rect -198 -144960 -94 -144761
rect 282 -144812 302 -140578
rect 366 -144812 386 -140578
rect 282 -144960 386 -144812
<< properties >>
string FIXED_BBOX -386 140550 94 144840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 64 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
