magic
tech sky130A
magscale 1 2
timestamp 1665169768
<< error_p >>
rect -87361 51620 -87301 56030
rect -87281 51620 -87221 56030
rect -86642 51620 -86582 56030
rect -86562 51620 -86502 56030
rect -85923 51620 -85863 56030
rect -85843 51620 -85783 56030
rect -85204 51620 -85144 56030
rect -85124 51620 -85064 56030
rect -84485 51620 -84425 56030
rect -84405 51620 -84345 56030
rect -83766 51620 -83706 56030
rect -83686 51620 -83626 56030
rect -83047 51620 -82987 56030
rect -82967 51620 -82907 56030
rect -82328 51620 -82268 56030
rect -82248 51620 -82188 56030
rect -81609 51620 -81549 56030
rect -81529 51620 -81469 56030
rect -80890 51620 -80830 56030
rect -80810 51620 -80750 56030
rect -80171 51620 -80111 56030
rect -80091 51620 -80031 56030
rect -79452 51620 -79392 56030
rect -79372 51620 -79312 56030
rect -78733 51620 -78673 56030
rect -78653 51620 -78593 56030
rect -78014 51620 -77954 56030
rect -77934 51620 -77874 56030
rect -77295 51620 -77260 56030
rect -68642 51620 -68582 56030
rect -68562 51620 -68502 56030
rect -67923 51620 -67863 56030
rect -67843 51620 -67783 56030
rect -67204 51620 -67144 56030
rect -67124 51620 -67064 56030
rect -66485 51620 -66425 56030
rect -66405 51620 -66345 56030
rect -65766 51620 -65706 56030
rect -65686 51620 -65626 56030
rect -65047 51620 -64987 56030
rect -64967 51620 -64907 56030
rect -64328 51620 -64268 56030
rect -64248 51620 -64188 56030
rect -63609 51620 -63549 56030
rect -63529 51620 -63469 56030
rect -62890 51620 -62830 56030
rect -62810 51620 -62750 56030
rect -62171 51620 -62111 56030
rect -62091 51620 -62031 56030
rect -61452 51620 -61392 56030
rect -61372 51620 -61312 56030
rect -60733 51620 -60673 56030
rect -60653 51620 -60593 56030
rect -60014 51620 -59954 56030
rect -59934 51620 -59874 56030
rect -59295 51620 -59260 56030
rect -43361 51620 -43301 56030
rect -43281 51620 -43221 56030
rect -42642 51620 -42582 56030
rect -42562 51620 -42502 56030
rect -41923 51620 -41863 56030
rect -41843 51620 -41783 56030
rect -87361 47110 -87301 51520
rect -87281 47110 -87221 51520
rect -86642 47110 -86582 51520
rect -86562 47110 -86502 51520
rect -85923 47110 -85863 51520
rect -85843 47110 -85783 51520
rect -85204 47110 -85144 51520
rect -85124 47110 -85064 51520
rect -84485 47110 -84425 51520
rect -84405 47110 -84345 51520
rect -83766 47110 -83706 51520
rect -83686 47110 -83626 51520
rect -83047 47110 -82987 51520
rect -82967 47110 -82907 51520
rect -82328 47110 -82268 51520
rect -82248 47110 -82188 51520
rect -81609 47110 -81549 51520
rect -81529 47110 -81469 51520
rect -80890 47110 -80830 51520
rect -80810 47110 -80750 51520
rect -80171 47110 -80111 51520
rect -80091 47110 -80031 51520
rect -79452 47110 -79392 51520
rect -79372 47110 -79312 51520
rect -78733 47110 -78673 51520
rect -78653 47110 -78593 51520
rect -78014 47110 -77954 51520
rect -77934 47110 -77874 51520
rect -77295 47110 -77260 51520
rect -68642 47110 -68582 51520
rect -68562 47110 -68502 51520
rect -67923 47110 -67863 51520
rect -67843 47110 -67783 51520
rect -67204 47110 -67144 51520
rect -67124 47110 -67064 51520
rect -66485 47110 -66425 51520
rect -66405 47110 -66345 51520
rect -65766 47110 -65706 51520
rect -65686 47110 -65626 51520
rect -65047 47110 -64987 51520
rect -64967 47110 -64907 51520
rect -64328 47110 -64268 51520
rect -64248 47110 -64188 51520
rect -63609 47110 -63549 51520
rect -63529 47110 -63469 51520
rect -62890 47110 -62830 51520
rect -62810 47110 -62750 51520
rect -62171 47110 -62111 51520
rect -62091 47110 -62031 51520
rect -61452 47110 -61392 51520
rect -61372 47110 -61312 51520
rect -60733 47110 -60673 51520
rect -60653 47110 -60593 51520
rect -60014 47110 -59954 51520
rect -59934 47110 -59874 51520
rect -59295 47110 -59260 51520
rect -43361 47110 -43301 51520
rect -43281 47110 -43221 51520
rect -42642 47110 -42582 51520
rect -42562 47110 -42502 51520
rect -41923 47110 -41863 51520
rect -41843 47110 -41783 51520
rect -87361 42600 -87301 47010
rect -87281 42600 -87221 47010
rect -86642 42600 -86582 47010
rect -86562 42600 -86502 47010
rect -85923 42600 -85863 47010
rect -85843 42600 -85783 47010
rect -85204 42600 -85144 47010
rect -85124 42600 -85064 47010
rect -84485 42600 -84425 47010
rect -84405 42600 -84345 47010
rect -83766 42600 -83706 47010
rect -83686 42600 -83626 47010
rect -83047 42600 -82987 47010
rect -82967 42600 -82907 47010
rect -82328 42600 -82268 47010
rect -82248 42600 -82188 47010
rect -81609 42600 -81549 47010
rect -81529 42600 -81469 47010
rect -80890 42600 -80830 47010
rect -80810 42600 -80750 47010
rect -80171 42600 -80111 47010
rect -80091 42600 -80031 47010
rect -79452 42600 -79392 47010
rect -79372 42600 -79312 47010
rect -78733 42600 -78673 47010
rect -78653 42600 -78593 47010
rect -78014 42600 -77954 47010
rect -77934 42600 -77874 47010
rect -77295 42600 -77260 47010
rect -68642 42600 -68582 47010
rect -68562 42600 -68502 47010
rect -67923 42600 -67863 47010
rect -67843 42600 -67783 47010
rect -67204 42600 -67144 47010
rect -67124 42600 -67064 47010
rect -66485 42600 -66425 47010
rect -66405 42600 -66345 47010
rect -65766 42600 -65706 47010
rect -65686 42600 -65626 47010
rect -65047 42600 -64987 47010
rect -64967 42600 -64907 47010
rect -64328 42600 -64268 47010
rect -64248 42600 -64188 47010
rect -63609 42600 -63549 47010
rect -63529 42600 -63469 47010
rect -62890 42600 -62830 47010
rect -62810 42600 -62750 47010
rect -62171 42600 -62111 47010
rect -62091 42600 -62031 47010
rect -61452 42600 -61392 47010
rect -61372 42600 -61312 47010
rect -60733 42600 -60673 47010
rect -60653 42600 -60593 47010
rect -60014 42600 -59954 47010
rect -59934 42600 -59874 47010
rect -59295 42600 -59260 47010
rect -43361 42600 -43301 47010
rect -43281 42600 -43221 47010
rect -42642 42600 -42582 47010
rect -42562 42600 -42502 47010
rect -41923 42600 -41863 47010
rect -41843 42600 -41783 47010
rect -87361 38090 -87301 42500
rect -87281 38090 -87221 42500
rect -86642 38090 -86582 42500
rect -86562 38090 -86502 42500
rect -85923 38090 -85863 42500
rect -85843 38090 -85783 42500
rect -85204 38090 -85144 42500
rect -85124 38090 -85064 42500
rect -84485 38090 -84425 42500
rect -84405 38090 -84345 42500
rect -83766 38090 -83706 42500
rect -83686 38090 -83626 42500
rect -83047 38090 -82987 42500
rect -82967 38090 -82907 42500
rect -82328 38090 -82268 42500
rect -82248 38090 -82188 42500
rect -81609 38090 -81549 42500
rect -81529 38090 -81469 42500
rect -80890 38090 -80830 42500
rect -80810 38090 -80750 42500
rect -80171 38090 -80111 42500
rect -80091 38090 -80031 42500
rect -79452 38090 -79392 42500
rect -79372 38090 -79312 42500
rect -78733 38090 -78673 42500
rect -78653 38090 -78593 42500
rect -78014 38090 -77954 42500
rect -77934 38090 -77874 42500
rect -77295 38090 -77260 42500
rect -68642 38090 -68582 42500
rect -68562 38090 -68502 42500
rect -67923 38090 -67863 42500
rect -67843 38090 -67783 42500
rect -67204 38090 -67144 42500
rect -67124 38090 -67064 42500
rect -66485 38090 -66425 42500
rect -66405 38090 -66345 42500
rect -65766 38090 -65706 42500
rect -65686 38090 -65626 42500
rect -65047 38090 -64987 42500
rect -64967 38090 -64907 42500
rect -64328 38090 -64268 42500
rect -64248 38090 -64188 42500
rect -63609 38090 -63549 42500
rect -63529 38090 -63469 42500
rect -62890 38090 -62830 42500
rect -62810 38090 -62750 42500
rect -62171 38090 -62111 42500
rect -62091 38090 -62031 42500
rect -61452 38090 -61392 42500
rect -61372 38090 -61312 42500
rect -60733 38090 -60673 42500
rect -60653 38090 -60593 42500
rect -60014 38090 -59954 42500
rect -59934 38090 -59874 42500
rect -59295 38090 -59260 42500
rect -43361 38090 -43301 42500
rect -43281 38090 -43221 42500
rect -42642 38090 -42582 42500
rect -42562 38090 -42502 42500
rect -41923 38090 -41863 42500
rect -41843 38090 -41783 42500
rect -87361 33580 -87301 37990
rect -87281 33580 -87221 37990
rect -86642 33580 -86582 37990
rect -86562 33580 -86502 37990
rect -85923 33580 -85863 37990
rect -85843 33580 -85783 37990
rect -85204 33580 -85144 37990
rect -85124 33580 -85064 37990
rect -84485 33580 -84425 37990
rect -84405 33580 -84345 37990
rect -83766 33580 -83706 37990
rect -83686 33580 -83626 37990
rect -83047 33580 -82987 37990
rect -82967 33580 -82907 37990
rect -82328 33580 -82268 37990
rect -82248 33580 -82188 37990
rect -81609 33580 -81549 37990
rect -81529 33580 -81469 37990
rect -80890 33580 -80830 37990
rect -80810 33580 -80750 37990
rect -80171 33580 -80111 37990
rect -80091 33580 -80031 37990
rect -79452 33580 -79392 37990
rect -79372 33580 -79312 37990
rect -78733 33580 -78673 37990
rect -78653 33580 -78593 37990
rect -78014 33580 -77954 37990
rect -77934 33580 -77874 37990
rect -77295 33580 -77260 37990
rect -68642 33580 -68582 37990
rect -68562 33580 -68502 37990
rect -67923 33580 -67863 37990
rect -67843 33580 -67783 37990
rect -67204 33580 -67144 37990
rect -67124 33580 -67064 37990
rect -66485 33580 -66425 37990
rect -66405 33580 -66345 37990
rect -65766 33580 -65706 37990
rect -65686 33580 -65626 37990
rect -65047 33580 -64987 37990
rect -64967 33580 -64907 37990
rect -64328 33580 -64268 37990
rect -64248 33580 -64188 37990
rect -63609 33580 -63549 37990
rect -63529 33580 -63469 37990
rect -62890 33580 -62830 37990
rect -62810 33580 -62750 37990
rect -62171 33580 -62111 37990
rect -62091 33580 -62031 37990
rect -61452 33580 -61392 37990
rect -61372 33580 -61312 37990
rect -60733 33580 -60673 37990
rect -60653 33580 -60593 37990
rect -60014 33580 -59954 37990
rect -59934 33580 -59874 37990
rect -59295 33580 -59260 37990
rect -43361 33580 -43301 37990
rect -43281 33580 -43221 37990
rect -42642 33580 -42582 37990
rect -42562 33580 -42502 37990
rect -41923 33580 -41863 37990
rect -41843 33580 -41783 37990
rect -87361 29070 -87301 33480
rect -87281 29070 -87221 33480
rect -86642 29070 -86582 33480
rect -86562 29070 -86502 33480
rect -85923 29070 -85863 33480
rect -85843 29070 -85783 33480
rect -85204 29070 -85144 33480
rect -85124 29070 -85064 33480
rect -84485 29070 -84425 33480
rect -84405 29070 -84345 33480
rect -83766 29070 -83706 33480
rect -83686 29070 -83626 33480
rect -83047 29070 -82987 33480
rect -82967 29070 -82907 33480
rect -82328 29070 -82268 33480
rect -82248 29070 -82188 33480
rect -81609 29070 -81549 33480
rect -81529 29070 -81469 33480
rect -80890 29070 -80830 33480
rect -80810 29070 -80750 33480
rect -80171 29070 -80111 33480
rect -80091 29070 -80031 33480
rect -79452 29070 -79392 33480
rect -79372 29070 -79312 33480
rect -78733 29070 -78673 33480
rect -78653 29070 -78593 33480
rect -78014 29070 -77954 33480
rect -77934 29070 -77874 33480
rect -77295 29070 -77260 33480
rect -68642 29070 -68582 33480
rect -68562 29070 -68502 33480
rect -67923 29070 -67863 33480
rect -67843 29070 -67783 33480
rect -67204 29070 -67144 33480
rect -67124 29070 -67064 33480
rect -66485 29070 -66425 33480
rect -66405 29070 -66345 33480
rect -65766 29070 -65706 33480
rect -65686 29070 -65626 33480
rect -65047 29070 -64987 33480
rect -64967 29070 -64907 33480
rect -64328 29070 -64268 33480
rect -64248 29070 -64188 33480
rect -63609 29070 -63549 33480
rect -63529 29070 -63469 33480
rect -62890 29070 -62830 33480
rect -62810 29070 -62750 33480
rect -62171 29070 -62111 33480
rect -62091 29070 -62031 33480
rect -61452 29070 -61392 33480
rect -61372 29070 -61312 33480
rect -60733 29070 -60673 33480
rect -60653 29070 -60593 33480
rect -60014 29070 -59954 33480
rect -59934 29070 -59874 33480
rect -59295 29070 -59260 33480
rect -43361 29070 -43301 33480
rect -43281 29070 -43221 33480
rect -42642 29070 -42582 33480
rect -42562 29070 -42502 33480
rect -41923 29070 -41863 33480
rect -41843 29070 -41783 33480
rect -87361 24560 -87301 28970
rect -87281 24560 -87221 28970
rect -86642 24560 -86582 28970
rect -86562 24560 -86502 28970
rect -85923 24560 -85863 28970
rect -85843 24560 -85783 28970
rect -85204 24560 -85144 28970
rect -85124 24560 -85064 28970
rect -84485 24560 -84425 28970
rect -84405 24560 -84345 28970
rect -83766 24560 -83706 28970
rect -83686 24560 -83626 28970
rect -83047 24560 -82987 28970
rect -82967 24560 -82907 28970
rect -82328 24560 -82268 28970
rect -82248 24560 -82188 28970
rect -81609 24560 -81549 28970
rect -81529 24560 -81469 28970
rect -80890 24560 -80830 28970
rect -80810 24560 -80750 28970
rect -80171 24560 -80111 28970
rect -80091 24560 -80031 28970
rect -79452 24560 -79392 28970
rect -79372 24560 -79312 28970
rect -78733 24560 -78673 28970
rect -78653 24560 -78593 28970
rect -78014 24560 -77954 28970
rect -77934 24560 -77874 28970
rect -77295 24560 -77260 28970
rect -68642 24560 -68582 28970
rect -68562 24560 -68502 28970
rect -67923 24560 -67863 28970
rect -67843 24560 -67783 28970
rect -67204 24560 -67144 28970
rect -67124 24560 -67064 28970
rect -66485 24560 -66425 28970
rect -66405 24560 -66345 28970
rect -65766 24560 -65706 28970
rect -65686 24560 -65626 28970
rect -65047 24560 -64987 28970
rect -64967 24560 -64907 28970
rect -64328 24560 -64268 28970
rect -64248 24560 -64188 28970
rect -63609 24560 -63549 28970
rect -63529 24560 -63469 28970
rect -62890 24560 -62830 28970
rect -62810 24560 -62750 28970
rect -62171 24560 -62111 28970
rect -62091 24560 -62031 28970
rect -61452 24560 -61392 28970
rect -61372 24560 -61312 28970
rect -60733 24560 -60673 28970
rect -60653 24560 -60593 28970
rect -60014 24560 -59954 28970
rect -59934 24560 -59874 28970
rect -59295 24560 -59260 28970
rect -43361 24560 -43301 28970
rect -43281 24560 -43221 28970
rect -42642 24560 -42582 28970
rect -42562 24560 -42502 28970
rect -41923 24560 -41863 28970
rect -41843 24560 -41783 28970
rect -87361 20050 -87301 24460
rect -87281 20050 -87221 24460
rect -86642 20050 -86582 24460
rect -86562 20050 -86502 24460
rect -85923 20050 -85863 24460
rect -85843 20050 -85783 24460
rect -85204 20050 -85144 24460
rect -85124 20050 -85064 24460
rect -84485 20050 -84425 24460
rect -84405 20050 -84345 24460
rect -83766 20050 -83706 24460
rect -83686 20050 -83626 24460
rect -83047 20050 -82987 24460
rect -82967 20050 -82907 24460
rect -82328 20050 -82268 24460
rect -82248 20050 -82188 24460
rect -81609 20050 -81549 24460
rect -81529 20050 -81469 24460
rect -80890 20050 -80830 24460
rect -80810 20050 -80750 24460
rect -80171 20050 -80111 24460
rect -80091 20050 -80031 24460
rect -79452 20050 -79392 24460
rect -79372 20050 -79312 24460
rect -78733 20050 -78673 24460
rect -78653 20050 -78593 24460
rect -78014 20050 -77954 24460
rect -77934 20050 -77874 24460
rect -77295 20050 -77260 24460
rect -68642 20050 -68582 24460
rect -68562 20050 -68502 24460
rect -67923 20050 -67863 24460
rect -67843 20050 -67783 24460
rect -67204 20050 -67144 24460
rect -67124 20050 -67064 24460
rect -66485 20050 -66425 24460
rect -66405 20050 -66345 24460
rect -65766 20050 -65706 24460
rect -65686 20050 -65626 24460
rect -65047 20050 -64987 24460
rect -64967 20050 -64907 24460
rect -64328 20050 -64268 24460
rect -64248 20050 -64188 24460
rect -63609 20050 -63549 24460
rect -63529 20050 -63469 24460
rect -62890 20050 -62830 24460
rect -62810 20050 -62750 24460
rect -62171 20050 -62111 24460
rect -62091 20050 -62031 24460
rect -61452 20050 -61392 24460
rect -61372 20050 -61312 24460
rect -60733 20050 -60673 24460
rect -60653 20050 -60593 24460
rect -60014 20050 -59954 24460
rect -59934 20050 -59874 24460
rect -59295 20050 -59260 24460
rect -43361 20050 -43301 24460
rect -43281 20050 -43221 24460
rect -42642 20050 -42582 24460
rect -42562 20050 -42502 24460
rect -41923 20050 -41863 24460
rect -41843 20050 -41783 24460
rect -87361 13620 -87301 18030
rect -87281 13620 -87221 18030
rect -86642 13620 -86582 18030
rect -86562 13620 -86502 18030
rect -85923 13620 -85863 18030
rect -85843 13620 -85783 18030
rect -85204 13620 -85144 18030
rect -85124 13620 -85064 18030
rect -84485 13620 -84425 18030
rect -84405 13620 -84345 18030
rect -83766 13620 -83706 18030
rect -83686 13620 -83626 18030
rect -83047 13620 -82987 18030
rect -82967 13620 -82907 18030
rect -82328 13620 -82268 18030
rect -82248 13620 -82188 18030
rect -81609 13620 -81549 18030
rect -81529 13620 -81469 18030
rect -80890 13620 -80830 18030
rect -80810 13620 -80750 18030
rect -80171 13620 -80111 18030
rect -80091 13620 -80031 18030
rect -79452 13620 -79392 18030
rect -79372 13620 -79312 18030
rect -78733 13620 -78673 18030
rect -78653 13620 -78593 18030
rect -78014 13620 -77954 18030
rect -77934 13620 -77874 18030
rect -77295 13620 -77260 18030
rect -68642 13620 -68582 18030
rect -68562 13620 -68502 18030
rect -67923 13620 -67863 18030
rect -67843 13620 -67783 18030
rect -67204 13620 -67144 18030
rect -67124 13620 -67064 18030
rect -66485 13620 -66425 18030
rect -66405 13620 -66345 18030
rect -65766 13620 -65706 18030
rect -65686 13620 -65626 18030
rect -65047 13620 -64987 18030
rect -64967 13620 -64907 18030
rect -64328 13620 -64268 18030
rect -64248 13620 -64188 18030
rect -63609 13620 -63549 18030
rect -63529 13620 -63469 18030
rect -62890 13620 -62830 18030
rect -62810 13620 -62750 18030
rect -62171 13620 -62111 18030
rect -62091 13620 -62031 18030
rect -61452 13620 -61392 18030
rect -61372 13620 -61312 18030
rect -60733 13620 -60673 18030
rect -60653 13620 -60593 18030
rect -60014 13620 -59954 18030
rect -59934 13620 -59874 18030
rect -59295 13620 -59260 18030
rect -43361 13620 -43301 18030
rect -43281 13620 -43221 18030
rect -42642 13620 -42582 18030
rect -42562 13620 -42502 18030
rect -41923 13620 -41863 18030
rect -41843 13620 -41783 18030
rect -87361 9110 -87301 13520
rect -87281 9110 -87221 13520
rect -86642 9110 -86582 13520
rect -86562 9110 -86502 13520
rect -85923 9110 -85863 13520
rect -85843 9110 -85783 13520
rect -85204 9110 -85144 13520
rect -85124 9110 -85064 13520
rect -84485 9110 -84425 13520
rect -84405 9110 -84345 13520
rect -83766 9110 -83706 13520
rect -83686 9110 -83626 13520
rect -83047 9110 -82987 13520
rect -82967 9110 -82907 13520
rect -82328 9110 -82268 13520
rect -82248 9110 -82188 13520
rect -81609 9110 -81549 13520
rect -81529 9110 -81469 13520
rect -80890 9110 -80830 13520
rect -80810 9110 -80750 13520
rect -80171 9110 -80111 13520
rect -80091 9110 -80031 13520
rect -79452 9110 -79392 13520
rect -79372 9110 -79312 13520
rect -78733 9110 -78673 13520
rect -78653 9110 -78593 13520
rect -78014 9110 -77954 13520
rect -77934 9110 -77874 13520
rect -77295 9110 -77260 13520
rect -68642 9110 -68582 13520
rect -68562 9110 -68502 13520
rect -67923 9110 -67863 13520
rect -67843 9110 -67783 13520
rect -67204 9110 -67144 13520
rect -67124 9110 -67064 13520
rect -66485 9110 -66425 13520
rect -66405 9110 -66345 13520
rect -65766 9110 -65706 13520
rect -65686 9110 -65626 13520
rect -65047 9110 -64987 13520
rect -64967 9110 -64907 13520
rect -64328 9110 -64268 13520
rect -64248 9110 -64188 13520
rect -63609 9110 -63549 13520
rect -63529 9110 -63469 13520
rect -62890 9110 -62830 13520
rect -62810 9110 -62750 13520
rect -62171 9110 -62111 13520
rect -62091 9110 -62031 13520
rect -61452 9110 -61392 13520
rect -61372 9110 -61312 13520
rect -60733 9110 -60673 13520
rect -60653 9110 -60593 13520
rect -60014 9110 -59954 13520
rect -59934 9110 -59874 13520
rect -59295 9110 -59260 13520
rect -43361 9110 -43301 13520
rect -43281 9110 -43221 13520
rect -42642 9110 -42582 13520
rect -42562 9110 -42502 13520
rect -41923 9110 -41863 13520
rect -41843 9110 -41783 13520
rect -87361 4600 -87301 9010
rect -87281 4600 -87221 9010
rect -86642 4600 -86582 9010
rect -86562 4600 -86502 9010
rect -85923 4600 -85863 9010
rect -85843 4600 -85783 9010
rect -85204 4600 -85144 9010
rect -85124 4600 -85064 9010
rect -84485 4600 -84425 9010
rect -84405 4600 -84345 9010
rect -83766 4600 -83706 9010
rect -83686 4600 -83626 9010
rect -83047 4600 -82987 9010
rect -82967 4600 -82907 9010
rect -82328 4600 -82268 9010
rect -82248 4600 -82188 9010
rect -81609 4600 -81549 9010
rect -81529 4600 -81469 9010
rect -80890 4600 -80830 9010
rect -80810 4600 -80750 9010
rect -80171 4600 -80111 9010
rect -80091 4600 -80031 9010
rect -79452 4600 -79392 9010
rect -79372 4600 -79312 9010
rect -78733 4600 -78673 9010
rect -78653 4600 -78593 9010
rect -78014 4600 -77954 9010
rect -77934 4600 -77874 9010
rect -77295 4600 -77260 9010
rect -68642 4600 -68582 9010
rect -68562 4600 -68502 9010
rect -67923 4600 -67863 9010
rect -67843 4600 -67783 9010
rect -67204 4600 -67144 9010
rect -67124 4600 -67064 9010
rect -66485 4600 -66425 9010
rect -66405 4600 -66345 9010
rect -65766 4600 -65706 9010
rect -65686 4600 -65626 9010
rect -65047 4600 -64987 9010
rect -64967 4600 -64907 9010
rect -64328 4600 -64268 9010
rect -64248 4600 -64188 9010
rect -63609 4600 -63549 9010
rect -63529 4600 -63469 9010
rect -62890 4600 -62830 9010
rect -62810 4600 -62750 9010
rect -62171 4600 -62111 9010
rect -62091 4600 -62031 9010
rect -61452 4600 -61392 9010
rect -61372 4600 -61312 9010
rect -60733 4600 -60673 9010
rect -60653 4600 -60593 9010
rect -60014 4600 -59954 9010
rect -59934 4600 -59874 9010
rect -59295 4600 -59260 9010
rect -43361 4600 -43301 9010
rect -43281 4600 -43221 9010
rect -42642 4600 -42582 9010
rect -42562 4600 -42502 9010
rect -41923 4600 -41863 9010
rect -41843 4600 -41783 9010
rect -87361 90 -87301 4500
rect -87281 90 -87221 4500
rect -86642 90 -86582 4500
rect -86562 90 -86502 4500
rect -85923 90 -85863 4500
rect -85843 90 -85783 4500
rect -85204 90 -85144 4500
rect -85124 90 -85064 4500
rect -84485 90 -84425 4500
rect -84405 90 -84345 4500
rect -83766 90 -83706 4500
rect -83686 90 -83626 4500
rect -83047 90 -82987 4500
rect -82967 90 -82907 4500
rect -82328 90 -82268 4500
rect -82248 90 -82188 4500
rect -81609 90 -81549 4500
rect -81529 90 -81469 4500
rect -80890 90 -80830 4500
rect -80810 90 -80750 4500
rect -80171 90 -80111 4500
rect -80091 90 -80031 4500
rect -79452 90 -79392 4500
rect -79372 90 -79312 4500
rect -78733 90 -78673 4500
rect -78653 90 -78593 4500
rect -78014 90 -77954 4500
rect -77934 90 -77874 4500
rect -77295 90 -77260 4500
rect -68642 90 -68582 4500
rect -68562 90 -68502 4500
rect -67923 90 -67863 4500
rect -67843 90 -67783 4500
rect -67204 90 -67144 4500
rect -67124 90 -67064 4500
rect -66485 90 -66425 4500
rect -66405 90 -66345 4500
rect -65766 90 -65706 4500
rect -65686 90 -65626 4500
rect -65047 90 -64987 4500
rect -64967 90 -64907 4500
rect -64328 90 -64268 4500
rect -64248 90 -64188 4500
rect -63609 90 -63549 4500
rect -63529 90 -63469 4500
rect -62890 90 -62830 4500
rect -62810 90 -62750 4500
rect -62171 90 -62111 4500
rect -62091 90 -62031 4500
rect -61452 90 -61392 4500
rect -61372 90 -61312 4500
rect -60733 90 -60673 4500
rect -60653 90 -60593 4500
rect -60014 90 -59954 4500
rect -59934 90 -59874 4500
rect -59295 90 -59260 4500
rect -43361 90 -43301 4500
rect -43281 90 -43221 4500
rect -42642 90 -42582 4500
rect -42562 90 -42502 4500
rect -41923 90 -41863 4500
rect -41843 90 -41783 4500
rect -87361 -4420 -87301 -10
rect -87281 -4420 -87221 -10
rect -86642 -4420 -86582 -10
rect -86562 -4420 -86502 -10
rect -85923 -4420 -85863 -10
rect -85843 -4420 -85783 -10
rect -85204 -4420 -85144 -10
rect -85124 -4420 -85064 -10
rect -84485 -4420 -84425 -10
rect -84405 -4420 -84345 -10
rect -83766 -4420 -83706 -10
rect -83686 -4420 -83626 -10
rect -83047 -4420 -82987 -10
rect -82967 -4420 -82907 -10
rect -82328 -4420 -82268 -10
rect -82248 -4420 -82188 -10
rect -81609 -4420 -81549 -10
rect -81529 -4420 -81469 -10
rect -80890 -4420 -80830 -10
rect -80810 -4420 -80750 -10
rect -80171 -4420 -80111 -10
rect -80091 -4420 -80031 -10
rect -79452 -4420 -79392 -10
rect -79372 -4420 -79312 -10
rect -78733 -4420 -78673 -10
rect -78653 -4420 -78593 -10
rect -78014 -4420 -77954 -10
rect -77934 -4420 -77874 -10
rect -77295 -4420 -77260 -10
rect -75256 -4420 -75221 -10
rect -74642 -4420 -74582 -10
rect -74562 -4420 -74502 -10
rect -73923 -4420 -73863 -10
rect -73843 -4420 -73783 -10
rect -73204 -4420 -73144 -10
rect -73124 -4420 -73064 -10
rect -68642 -4420 -68582 -10
rect -68562 -4420 -68502 -10
rect -67923 -4420 -67863 -10
rect -67843 -4420 -67783 -10
rect -67204 -4420 -67144 -10
rect -67124 -4420 -67064 -10
rect -66485 -4420 -66425 -10
rect -66405 -4420 -66345 -10
rect -65766 -4420 -65706 -10
rect -65686 -4420 -65626 -10
rect -65047 -4420 -64987 -10
rect -64967 -4420 -64907 -10
rect -64328 -4420 -64268 -10
rect -64248 -4420 -64188 -10
rect -63609 -4420 -63549 -10
rect -63529 -4420 -63469 -10
rect -62890 -4420 -62830 -10
rect -62810 -4420 -62750 -10
rect -62171 -4420 -62111 -10
rect -62091 -4420 -62031 -10
rect -61452 -4420 -61392 -10
rect -61372 -4420 -61312 -10
rect -60733 -4420 -60673 -10
rect -60653 -4420 -60593 -10
rect -60014 -4420 -59954 -10
rect -59934 -4420 -59874 -10
rect -59295 -4420 -59260 -10
rect -43361 -4420 -43301 -10
rect -43281 -4420 -43221 -10
rect -42642 -4420 -42582 -10
rect -42562 -4420 -42502 -10
rect -41923 -4420 -41863 -10
rect -41843 -4420 -41783 -10
rect -87361 -8930 -87301 -4520
rect -87281 -8930 -87221 -4520
rect -86642 -8930 -86582 -4520
rect -86562 -8930 -86502 -4520
rect -85923 -8930 -85863 -4520
rect -85843 -8930 -85783 -4520
rect -85204 -8930 -85144 -4520
rect -85124 -8930 -85064 -4520
rect -84485 -8930 -84425 -4520
rect -84405 -8930 -84345 -4520
rect -83766 -8930 -83706 -4520
rect -83686 -8930 -83626 -4520
rect -83047 -8930 -82987 -4520
rect -82967 -8930 -82907 -4520
rect -82328 -8930 -82268 -4520
rect -82248 -8930 -82188 -4520
rect -81609 -8930 -81549 -4520
rect -81529 -8930 -81469 -4520
rect -80890 -8930 -80830 -4520
rect -80810 -8930 -80750 -4520
rect -80171 -8930 -80111 -4520
rect -80091 -8930 -80031 -4520
rect -79452 -8930 -79392 -4520
rect -79372 -8930 -79312 -4520
rect -78733 -8930 -78673 -4520
rect -78653 -8930 -78593 -4520
rect -78014 -8930 -77954 -4520
rect -77934 -8930 -77874 -4520
rect -77295 -8930 -77260 -4520
rect -75256 -8930 -75221 -4520
rect -74642 -8930 -74582 -4520
rect -74562 -8930 -74502 -4520
rect -73923 -8930 -73863 -4520
rect -73843 -8930 -73783 -4520
rect -73204 -8930 -73144 -4520
rect -73124 -8930 -73064 -4520
rect -68642 -8930 -68582 -4520
rect -68562 -8930 -68502 -4520
rect -67923 -8930 -67863 -4520
rect -67843 -8930 -67783 -4520
rect -67204 -8930 -67144 -4520
rect -67124 -8930 -67064 -4520
rect -66485 -8930 -66425 -4520
rect -66405 -8930 -66345 -4520
rect -65766 -8930 -65706 -4520
rect -65686 -8930 -65626 -4520
rect -65047 -8930 -64987 -4520
rect -64967 -8930 -64907 -4520
rect -64328 -8930 -64268 -4520
rect -64248 -8930 -64188 -4520
rect -63609 -8930 -63549 -4520
rect -63529 -8930 -63469 -4520
rect -62890 -8930 -62830 -4520
rect -62810 -8930 -62750 -4520
rect -62171 -8930 -62111 -4520
rect -62091 -8930 -62031 -4520
rect -61452 -8930 -61392 -4520
rect -61372 -8930 -61312 -4520
rect -60733 -8930 -60673 -4520
rect -60653 -8930 -60593 -4520
rect -60014 -8930 -59954 -4520
rect -59934 -8930 -59874 -4520
rect -59295 -8930 -59260 -4520
rect -43361 -8930 -43301 -4520
rect -43281 -8930 -43221 -4520
rect -42642 -8930 -42582 -4520
rect -42562 -8930 -42502 -4520
rect -41923 -8930 -41863 -4520
rect -41843 -8930 -41783 -4520
rect -87361 -13440 -87301 -9030
rect -87281 -13440 -87221 -9030
rect -86642 -13440 -86582 -9030
rect -86562 -13440 -86502 -9030
rect -85923 -13440 -85863 -9030
rect -85843 -13440 -85783 -9030
rect -85204 -13440 -85144 -9030
rect -85124 -13440 -85064 -9030
rect -84485 -13440 -84425 -9030
rect -84405 -13440 -84345 -9030
rect -83766 -13440 -83706 -9030
rect -83686 -13440 -83626 -9030
rect -83047 -13440 -82987 -9030
rect -82967 -13440 -82907 -9030
rect -82328 -13440 -82268 -9030
rect -82248 -13440 -82188 -9030
rect -81609 -13440 -81549 -9030
rect -81529 -13440 -81469 -9030
rect -80890 -13440 -80830 -9030
rect -80810 -13440 -80750 -9030
rect -80171 -13440 -80111 -9030
rect -80091 -13440 -80031 -9030
rect -79452 -13440 -79392 -9030
rect -79372 -13440 -79312 -9030
rect -78733 -13440 -78673 -9030
rect -78653 -13440 -78593 -9030
rect -78014 -13440 -77954 -9030
rect -77934 -13440 -77874 -9030
rect -77295 -13440 -77260 -9030
rect -75256 -13440 -75221 -9030
rect -74642 -13440 -74582 -9030
rect -74562 -13440 -74502 -9030
rect -73923 -13440 -73863 -9030
rect -73843 -13440 -73783 -9030
rect -73204 -13440 -73144 -9030
rect -73124 -13440 -73064 -9030
rect -68642 -13440 -68582 -9030
rect -68562 -13440 -68502 -9030
rect -67923 -13440 -67863 -9030
rect -67843 -13440 -67783 -9030
rect -67204 -13440 -67144 -9030
rect -67124 -13440 -67064 -9030
rect -66485 -13440 -66425 -9030
rect -66405 -13440 -66345 -9030
rect -65766 -13440 -65706 -9030
rect -65686 -13440 -65626 -9030
rect -65047 -13440 -64987 -9030
rect -64967 -13440 -64907 -9030
rect -64328 -13440 -64268 -9030
rect -64248 -13440 -64188 -9030
rect -63609 -13440 -63549 -9030
rect -63529 -13440 -63469 -9030
rect -62890 -13440 -62830 -9030
rect -62810 -13440 -62750 -9030
rect -62171 -13440 -62111 -9030
rect -62091 -13440 -62031 -9030
rect -61452 -13440 -61392 -9030
rect -61372 -13440 -61312 -9030
rect -60733 -13440 -60673 -9030
rect -60653 -13440 -60593 -9030
rect -60014 -13440 -59954 -9030
rect -59934 -13440 -59874 -9030
rect -59295 -13440 -59260 -9030
rect -43361 -13440 -43301 -9030
rect -43281 -13440 -43221 -9030
rect -42642 -13440 -42582 -9030
rect -42562 -13440 -42502 -9030
rect -41923 -13440 -41863 -9030
rect -41843 -13440 -41783 -9030
rect -87361 -17950 -87301 -13540
rect -87281 -17950 -87221 -13540
rect -86642 -17950 -86582 -13540
rect -86562 -17950 -86502 -13540
rect -85923 -17950 -85863 -13540
rect -85843 -17950 -85783 -13540
rect -85204 -17950 -85144 -13540
rect -85124 -17950 -85064 -13540
rect -84485 -17950 -84425 -13540
rect -84405 -17950 -84345 -13540
rect -83766 -17950 -83706 -13540
rect -83686 -17950 -83626 -13540
rect -83047 -17950 -82987 -13540
rect -82967 -17950 -82907 -13540
rect -82328 -17950 -82268 -13540
rect -82248 -17950 -82188 -13540
rect -81609 -17950 -81549 -13540
rect -81529 -17950 -81469 -13540
rect -80890 -17950 -80830 -13540
rect -80810 -17950 -80750 -13540
rect -80171 -17950 -80111 -13540
rect -80091 -17950 -80031 -13540
rect -79452 -17950 -79392 -13540
rect -79372 -17950 -79312 -13540
rect -78733 -17950 -78673 -13540
rect -78653 -17950 -78593 -13540
rect -78014 -17950 -77954 -13540
rect -77934 -17950 -77874 -13540
rect -77295 -17950 -77260 -13540
rect -75256 -17950 -75221 -13540
rect -74642 -17950 -74582 -13540
rect -74562 -17950 -74502 -13540
rect -73923 -17950 -73863 -13540
rect -73843 -17950 -73783 -13540
rect -73204 -17950 -73144 -13540
rect -73124 -17950 -73064 -13540
rect -68642 -17950 -68582 -13540
rect -68562 -17950 -68502 -13540
rect -67923 -17950 -67863 -13540
rect -67843 -17950 -67783 -13540
rect -67204 -17950 -67144 -13540
rect -67124 -17950 -67064 -13540
rect -66485 -17950 -66425 -13540
rect -66405 -17950 -66345 -13540
rect -65766 -17950 -65706 -13540
rect -65686 -17950 -65626 -13540
rect -65047 -17950 -64987 -13540
rect -64967 -17950 -64907 -13540
rect -64328 -17950 -64268 -13540
rect -64248 -17950 -64188 -13540
rect -63609 -17950 -63549 -13540
rect -63529 -17950 -63469 -13540
rect -62890 -17950 -62830 -13540
rect -62810 -17950 -62750 -13540
rect -62171 -17950 -62111 -13540
rect -62091 -17950 -62031 -13540
rect -61452 -17950 -61392 -13540
rect -61372 -17950 -61312 -13540
rect -60733 -17950 -60673 -13540
rect -60653 -17950 -60593 -13540
rect -60014 -17950 -59954 -13540
rect -59934 -17950 -59874 -13540
rect -59295 -17950 -59260 -13540
rect -43361 -17950 -43301 -13540
rect -43281 -17950 -43221 -13540
rect -42642 -17950 -42582 -13540
rect -42562 -17950 -42502 -13540
rect -41923 -17950 -41863 -13540
rect -41843 -17950 -41783 -13540
<< error_s >>
rect -77260 51620 -77235 56030
rect -77215 51620 -77155 56030
rect -75361 51620 -75301 56030
rect -75281 51620 -75221 56030
rect -74642 51620 -74582 56030
rect -74562 51620 -74502 56030
rect -73923 51620 -73863 56030
rect -73843 51620 -73783 56030
rect -73204 51620 -73144 56030
rect -73124 51620 -73064 56030
rect -72485 51620 -72425 56030
rect -72405 51620 -72345 56030
rect -71766 51620 -71706 56030
rect -71686 51620 -71626 56030
rect -71047 51620 -70987 56030
rect -70967 51620 -70907 56030
rect -69361 51620 -69301 56030
rect -69281 51620 -69221 56030
rect -59260 51620 -59235 56030
rect -59215 51620 -59155 56030
rect -57361 51620 -57301 56030
rect -57281 51620 -57221 56030
rect -56642 51620 -56582 56030
rect -56562 51620 -56502 56030
rect -55923 51620 -55863 56030
rect -55843 51620 -55783 56030
rect -55204 51620 -55144 56030
rect -55124 51620 -55064 56030
rect -54485 51620 -54425 56030
rect -54405 51620 -54345 56030
rect -53766 51620 -53706 56030
rect -53686 51620 -53626 56030
rect -53047 51620 -52987 56030
rect -52967 51620 -52907 56030
rect -39361 51620 -39301 56030
rect -39281 51620 -39221 56030
rect -38642 51620 -38582 56030
rect -38562 51620 -38502 56030
rect -37923 51620 -37863 56030
rect -37843 51620 -37783 56030
rect -35361 51620 -35301 56030
rect -35281 51620 -35221 56030
rect -33361 51620 -33301 56030
rect -33281 51620 -33221 56030
rect -77260 47110 -77235 51520
rect -77215 47110 -77155 51520
rect -75361 47110 -75301 51520
rect -75281 47110 -75221 51520
rect -74642 47110 -74582 51520
rect -74562 47110 -74502 51520
rect -73923 47110 -73863 51520
rect -73843 47110 -73783 51520
rect -73204 47110 -73144 51520
rect -73124 47110 -73064 51520
rect -72485 47110 -72425 51520
rect -72405 47110 -72345 51520
rect -71766 47110 -71706 51520
rect -71686 47110 -71626 51520
rect -71047 47110 -70987 51520
rect -70967 47110 -70907 51520
rect -69361 47110 -69301 51520
rect -69281 47110 -69221 51520
rect -59260 47110 -59235 51520
rect -59215 47110 -59155 51520
rect -57361 47110 -57301 51520
rect -57281 47110 -57221 51520
rect -56642 47110 -56582 51520
rect -56562 47110 -56502 51520
rect -55923 47110 -55863 51520
rect -55843 47110 -55783 51520
rect -55204 47110 -55144 51520
rect -55124 47110 -55064 51520
rect -54485 47110 -54425 51520
rect -54405 47110 -54345 51520
rect -53766 47110 -53706 51520
rect -53686 47110 -53626 51520
rect -53047 47110 -52987 51520
rect -52967 47110 -52907 51520
rect -39361 47110 -39301 51520
rect -39281 47110 -39221 51520
rect -38642 47110 -38582 51520
rect -38562 47110 -38502 51520
rect -37923 47110 -37863 51520
rect -37843 47110 -37783 51520
rect -35361 47110 -35301 51520
rect -35281 47110 -35221 51520
rect -33361 47110 -33301 51520
rect -33281 47110 -33221 51520
rect -77260 42600 -77235 47010
rect -77215 42600 -77155 47010
rect -75361 42600 -75301 47010
rect -75281 42600 -75221 47010
rect -74642 42600 -74582 47010
rect -74562 42600 -74502 47010
rect -73923 42600 -73863 47010
rect -73843 42600 -73783 47010
rect -73204 42600 -73144 47010
rect -73124 42600 -73064 47010
rect -72485 42600 -72425 47010
rect -72405 42600 -72345 47010
rect -71766 42600 -71706 47010
rect -71686 42600 -71626 47010
rect -71047 42600 -70987 47010
rect -70967 42600 -70907 47010
rect -69361 42600 -69301 47010
rect -69281 42600 -69221 47010
rect -59260 42600 -59235 47010
rect -59215 42600 -59155 47010
rect -57361 42600 -57301 47010
rect -57281 42600 -57221 47010
rect -56642 42600 -56582 47010
rect -56562 42600 -56502 47010
rect -55923 42600 -55863 47010
rect -55843 42600 -55783 47010
rect -55204 42600 -55144 47010
rect -55124 42600 -55064 47010
rect -54485 42600 -54425 47010
rect -54405 42600 -54345 47010
rect -53766 42600 -53706 47010
rect -53686 42600 -53626 47010
rect -53047 42600 -52987 47010
rect -52967 42600 -52907 47010
rect -39361 42600 -39301 47010
rect -39281 42600 -39221 47010
rect -38642 42600 -38582 47010
rect -38562 42600 -38502 47010
rect -37923 42600 -37863 47010
rect -37843 42600 -37783 47010
rect -35361 42600 -35301 47010
rect -35281 42600 -35221 47010
rect -33361 42600 -33301 47010
rect -33281 42600 -33221 47010
rect -77260 38090 -77235 42500
rect -77215 38090 -77155 42500
rect -75361 38090 -75301 42500
rect -75281 38090 -75221 42500
rect -74642 38090 -74582 42500
rect -74562 38090 -74502 42500
rect -73923 38090 -73863 42500
rect -73843 38090 -73783 42500
rect -73204 38090 -73144 42500
rect -73124 38090 -73064 42500
rect -72485 38090 -72425 42500
rect -72405 38090 -72345 42500
rect -71766 38090 -71706 42500
rect -71686 38090 -71626 42500
rect -71047 38090 -70987 42500
rect -70967 38090 -70907 42500
rect -69361 38090 -69301 42500
rect -69281 38090 -69221 42500
rect -59260 38090 -59235 42500
rect -59215 38090 -59155 42500
rect -57361 38090 -57301 42500
rect -57281 38090 -57221 42500
rect -56642 38090 -56582 42500
rect -56562 38090 -56502 42500
rect -55923 38090 -55863 42500
rect -55843 38090 -55783 42500
rect -55204 38090 -55144 42500
rect -55124 38090 -55064 42500
rect -54485 38090 -54425 42500
rect -54405 38090 -54345 42500
rect -53766 38090 -53706 42500
rect -53686 38090 -53626 42500
rect -53047 38090 -52987 42500
rect -52967 38090 -52907 42500
rect -39361 38090 -39301 42500
rect -39281 38090 -39221 42500
rect -38642 38090 -38582 42500
rect -38562 38090 -38502 42500
rect -37923 38090 -37863 42500
rect -37843 38090 -37783 42500
rect -35361 38090 -35301 42500
rect -35281 38090 -35221 42500
rect -33361 38090 -33301 42500
rect -33281 38090 -33221 42500
rect -77260 33580 -77235 37990
rect -77215 33580 -77155 37990
rect -75361 33580 -75301 37990
rect -75281 33580 -75221 37990
rect -74642 33580 -74582 37990
rect -74562 33580 -74502 37990
rect -73923 33580 -73863 37990
rect -73843 33580 -73783 37990
rect -73204 33580 -73144 37990
rect -73124 33580 -73064 37990
rect -72485 33580 -72425 37990
rect -72405 33580 -72345 37990
rect -71766 33580 -71706 37990
rect -71686 33580 -71626 37990
rect -71047 33580 -70987 37990
rect -70967 33580 -70907 37990
rect -69361 33580 -69301 37990
rect -69281 33580 -69221 37990
rect -59260 33580 -59235 37990
rect -59215 33580 -59155 37990
rect -57361 33580 -57301 37990
rect -57281 33580 -57221 37990
rect -56642 33580 -56582 37990
rect -56562 33580 -56502 37990
rect -55923 33580 -55863 37990
rect -55843 33580 -55783 37990
rect -55204 33580 -55144 37990
rect -55124 33580 -55064 37990
rect -54485 33580 -54425 37990
rect -54405 33580 -54345 37990
rect -53766 33580 -53706 37990
rect -53686 33580 -53626 37990
rect -53047 33580 -52987 37990
rect -52967 33580 -52907 37990
rect -39361 33580 -39301 37990
rect -39281 33580 -39221 37990
rect -38642 33580 -38582 37990
rect -38562 33580 -38502 37990
rect -37923 33580 -37863 37990
rect -37843 33580 -37783 37990
rect -35361 33580 -35301 37990
rect -35281 33580 -35221 37990
rect -33361 33580 -33301 37990
rect -33281 33580 -33221 37990
rect -77260 29070 -77235 33480
rect -77215 29070 -77155 33480
rect -75361 29070 -75301 33480
rect -75281 29070 -75221 33480
rect -74642 29070 -74582 33480
rect -74562 29070 -74502 33480
rect -73923 29070 -73863 33480
rect -73843 29070 -73783 33480
rect -73204 29070 -73144 33480
rect -73124 29070 -73064 33480
rect -72485 29070 -72425 33480
rect -72405 29070 -72345 33480
rect -71766 29070 -71706 33480
rect -71686 29070 -71626 33480
rect -71047 29070 -70987 33480
rect -70967 29070 -70907 33480
rect -69361 29070 -69301 33480
rect -69281 29070 -69221 33480
rect -59260 29070 -59235 33480
rect -59215 29070 -59155 33480
rect -57361 29070 -57301 33480
rect -57281 29070 -57221 33480
rect -56642 29070 -56582 33480
rect -56562 29070 -56502 33480
rect -55923 29070 -55863 33480
rect -55843 29070 -55783 33480
rect -55204 29070 -55144 33480
rect -55124 29070 -55064 33480
rect -54485 29070 -54425 33480
rect -54405 29070 -54345 33480
rect -53766 29070 -53706 33480
rect -53686 29070 -53626 33480
rect -53047 29070 -52987 33480
rect -52967 29070 -52907 33480
rect -39361 29070 -39301 33480
rect -39281 29070 -39221 33480
rect -38642 29070 -38582 33480
rect -38562 29070 -38502 33480
rect -37923 29070 -37863 33480
rect -37843 29070 -37783 33480
rect -35361 29070 -35301 33480
rect -35281 29070 -35221 33480
rect -33361 29070 -33301 33480
rect -33281 29070 -33221 33480
rect -77260 24560 -77235 28970
rect -77215 24560 -77155 28970
rect -75361 24560 -75301 28970
rect -75281 24560 -75221 28970
rect -74642 24560 -74582 28970
rect -74562 24560 -74502 28970
rect -73923 24560 -73863 28970
rect -73843 24560 -73783 28970
rect -73204 24560 -73144 28970
rect -73124 24560 -73064 28970
rect -72485 24560 -72425 28970
rect -72405 24560 -72345 28970
rect -71766 24560 -71706 28970
rect -71686 24560 -71626 28970
rect -71047 24560 -70987 28970
rect -70967 24560 -70907 28970
rect -69361 24560 -69301 28970
rect -69281 24560 -69221 28970
rect -59260 24560 -59235 28970
rect -59215 24560 -59155 28970
rect -57361 24560 -57301 28970
rect -57281 24560 -57221 28970
rect -56642 24560 -56582 28970
rect -56562 24560 -56502 28970
rect -55923 24560 -55863 28970
rect -55843 24560 -55783 28970
rect -55204 24560 -55144 28970
rect -55124 24560 -55064 28970
rect -54485 24560 -54425 28970
rect -54405 24560 -54345 28970
rect -53766 24560 -53706 28970
rect -53686 24560 -53626 28970
rect -53047 24560 -52987 28970
rect -52967 24560 -52907 28970
rect -39361 24560 -39301 28970
rect -39281 24560 -39221 28970
rect -38642 24560 -38582 28970
rect -38562 24560 -38502 28970
rect -37923 24560 -37863 28970
rect -37843 24560 -37783 28970
rect -35361 24560 -35301 28970
rect -35281 24560 -35221 28970
rect -33361 24560 -33301 28970
rect -33281 24560 -33221 28970
rect -77260 20050 -77235 24460
rect -77215 20050 -77155 24460
rect -75361 20050 -75301 24460
rect -75281 20050 -75221 24460
rect -74642 20050 -74582 24460
rect -74562 20050 -74502 24460
rect -73923 20050 -73863 24460
rect -73843 20050 -73783 24460
rect -73204 20050 -73144 24460
rect -73124 20050 -73064 24460
rect -72485 20050 -72425 24460
rect -72405 20050 -72345 24460
rect -71766 20050 -71706 24460
rect -71686 20050 -71626 24460
rect -71047 20050 -70987 24460
rect -70967 20050 -70907 24460
rect -69361 20050 -69301 24460
rect -69281 20050 -69221 24460
rect -59260 20050 -59235 24460
rect -59215 20050 -59155 24460
rect -57361 20050 -57301 24460
rect -57281 20050 -57221 24460
rect -56642 20050 -56582 24460
rect -56562 20050 -56502 24460
rect -55923 20050 -55863 24460
rect -55843 20050 -55783 24460
rect -55204 20050 -55144 24460
rect -55124 20050 -55064 24460
rect -54485 20050 -54425 24460
rect -54405 20050 -54345 24460
rect -53766 20050 -53706 24460
rect -53686 20050 -53626 24460
rect -53047 20050 -52987 24460
rect -52967 20050 -52907 24460
rect -39361 20050 -39301 24460
rect -39281 20050 -39221 24460
rect -38642 20050 -38582 24460
rect -38562 20050 -38502 24460
rect -37923 20050 -37863 24460
rect -37843 20050 -37783 24460
rect -35361 20050 -35301 24460
rect -35281 20050 -35221 24460
rect -33361 20050 -33301 24460
rect -33281 20050 -33221 24460
rect -77260 13620 -77235 18030
rect -77215 13620 -77155 18030
rect -75361 13620 -75301 18030
rect -75281 13620 -75221 18030
rect -74642 13620 -74582 18030
rect -74562 13620 -74502 18030
rect -73923 13620 -73863 18030
rect -73843 13620 -73783 18030
rect -73204 13620 -73144 18030
rect -73124 13620 -73064 18030
rect -72485 13620 -72425 18030
rect -72405 13620 -72345 18030
rect -71766 13620 -71706 18030
rect -71686 13620 -71626 18030
rect -71047 13620 -70987 18030
rect -70967 13620 -70907 18030
rect -69361 13620 -69301 18030
rect -69281 13620 -69221 18030
rect -59260 13620 -59235 18030
rect -59215 13620 -59155 18030
rect -57361 13620 -57301 18030
rect -57281 13620 -57221 18030
rect -56642 13620 -56582 18030
rect -56562 13620 -56502 18030
rect -55923 13620 -55863 18030
rect -55843 13620 -55783 18030
rect -55204 13620 -55144 18030
rect -55124 13620 -55064 18030
rect -54485 13620 -54425 18030
rect -54405 13620 -54345 18030
rect -53766 13620 -53706 18030
rect -53686 13620 -53626 18030
rect -53047 13620 -52987 18030
rect -52967 13620 -52907 18030
rect -39361 13620 -39301 18030
rect -39281 13620 -39221 18030
rect -38642 13620 -38582 18030
rect -38562 13620 -38502 18030
rect -37923 13620 -37863 18030
rect -37843 13620 -37783 18030
rect -35361 13620 -35301 18030
rect -35281 13620 -35221 18030
rect -33361 13620 -33301 18030
rect -33281 13620 -33221 18030
rect -77260 9110 -77235 13520
rect -77215 9110 -77155 13520
rect -75361 9110 -75301 13520
rect -75281 9110 -75221 13520
rect -74642 9110 -74582 13520
rect -74562 9110 -74502 13520
rect -73923 9110 -73863 13520
rect -73843 9110 -73783 13520
rect -73204 9110 -73144 13520
rect -73124 9110 -73064 13520
rect -72485 9110 -72425 13520
rect -72405 9110 -72345 13520
rect -71766 9110 -71706 13520
rect -71686 9110 -71626 13520
rect -71047 9110 -70987 13520
rect -70967 9110 -70907 13520
rect -69361 9110 -69301 13520
rect -69281 9110 -69221 13520
rect -59260 9110 -59235 13520
rect -59215 9110 -59155 13520
rect -57361 9110 -57301 13520
rect -57281 9110 -57221 13520
rect -56642 9110 -56582 13520
rect -56562 9110 -56502 13520
rect -55923 9110 -55863 13520
rect -55843 9110 -55783 13520
rect -55204 9110 -55144 13520
rect -55124 9110 -55064 13520
rect -54485 9110 -54425 13520
rect -54405 9110 -54345 13520
rect -53766 9110 -53706 13520
rect -53686 9110 -53626 13520
rect -53047 9110 -52987 13520
rect -52967 9110 -52907 13520
rect -39361 9110 -39301 13520
rect -39281 9110 -39221 13520
rect -38642 9110 -38582 13520
rect -38562 9110 -38502 13520
rect -37923 9110 -37863 13520
rect -37843 9110 -37783 13520
rect -35361 9110 -35301 13520
rect -35281 9110 -35221 13520
rect -33361 9110 -33301 13520
rect -33281 9110 -33221 13520
rect -77260 4600 -77235 9010
rect -77215 4600 -77155 9010
rect -75361 4600 -75301 9010
rect -75281 4600 -75221 9010
rect -74642 4600 -74582 9010
rect -74562 4600 -74502 9010
rect -73923 4600 -73863 9010
rect -73843 4600 -73783 9010
rect -73204 4600 -73144 9010
rect -73124 4600 -73064 9010
rect -72485 4600 -72425 9010
rect -72405 4600 -72345 9010
rect -71766 4600 -71706 9010
rect -71686 4600 -71626 9010
rect -71047 4600 -70987 9010
rect -70967 4600 -70907 9010
rect -69361 4600 -69301 9010
rect -69281 4600 -69221 9010
rect -59260 4600 -59235 9010
rect -59215 4600 -59155 9010
rect -57361 4600 -57301 9010
rect -57281 4600 -57221 9010
rect -56642 4600 -56582 9010
rect -56562 4600 -56502 9010
rect -55923 4600 -55863 9010
rect -55843 4600 -55783 9010
rect -55204 4600 -55144 9010
rect -55124 4600 -55064 9010
rect -54485 4600 -54425 9010
rect -54405 4600 -54345 9010
rect -53766 4600 -53706 9010
rect -53686 4600 -53626 9010
rect -53047 4600 -52987 9010
rect -52967 4600 -52907 9010
rect -39361 4600 -39301 9010
rect -39281 4600 -39221 9010
rect -38642 4600 -38582 9010
rect -38562 4600 -38502 9010
rect -37923 4600 -37863 9010
rect -37843 4600 -37783 9010
rect -35361 4600 -35301 9010
rect -35281 4600 -35221 9010
rect -33361 4600 -33301 9010
rect -33281 4600 -33221 9010
rect -77260 90 -77235 4500
rect -77215 90 -77155 4500
rect -75361 90 -75301 4500
rect -75281 90 -75221 4500
rect -74642 90 -74582 4500
rect -74562 90 -74502 4500
rect -73923 90 -73863 4500
rect -73843 90 -73783 4500
rect -73204 90 -73144 4500
rect -73124 90 -73064 4500
rect -72485 90 -72425 4500
rect -72405 90 -72345 4500
rect -71766 90 -71706 4500
rect -71686 90 -71626 4500
rect -71047 90 -70987 4500
rect -70967 90 -70907 4500
rect -69361 90 -69301 4500
rect -69281 90 -69221 4500
rect -59260 90 -59235 4500
rect -59215 90 -59155 4500
rect -57361 90 -57301 4500
rect -57281 90 -57221 4500
rect -56642 90 -56582 4500
rect -56562 90 -56502 4500
rect -55923 90 -55863 4500
rect -55843 90 -55783 4500
rect -55204 90 -55144 4500
rect -55124 90 -55064 4500
rect -54485 90 -54425 4500
rect -54405 90 -54345 4500
rect -53766 90 -53706 4500
rect -53686 90 -53626 4500
rect -53047 90 -52987 4500
rect -52967 90 -52907 4500
rect -39361 90 -39301 4500
rect -39281 90 -39221 4500
rect -38642 90 -38582 4500
rect -38562 90 -38502 4500
rect -37923 90 -37863 4500
rect -37843 90 -37783 4500
rect -35361 90 -35301 4500
rect -35281 90 -35221 4500
rect -33361 90 -33301 4500
rect -33281 90 -33221 4500
rect -77260 -4420 -77235 -10
rect -77215 -4420 -77155 -10
rect -75361 -4420 -75301 -10
rect -75281 -4420 -75256 -10
rect -71047 -4420 -70987 -10
rect -70967 -4420 -70907 -10
rect -69361 -4420 -69301 -10
rect -69281 -4420 -69221 -10
rect -59260 -4420 -59235 -10
rect -59215 -4420 -59155 -10
rect -57361 -4420 -57301 -10
rect -57281 -4420 -57221 -10
rect -56642 -4420 -56582 -10
rect -56562 -4420 -56502 -10
rect -55923 -4420 -55863 -10
rect -55843 -4420 -55783 -10
rect -55204 -4420 -55144 -10
rect -55124 -4420 -55064 -10
rect -54485 -4420 -54425 -10
rect -54405 -4420 -54345 -10
rect -53766 -4420 -53706 -10
rect -53686 -4420 -53626 -10
rect -53047 -4420 -52987 -10
rect -52967 -4420 -52907 -10
rect -39361 -4420 -39301 -10
rect -39281 -4420 -39221 -10
rect -38642 -4420 -38582 -10
rect -38562 -4420 -38502 -10
rect -37923 -4420 -37863 -10
rect -37843 -4420 -37783 -10
rect -35361 -4420 -35301 -10
rect -35281 -4420 -35221 -10
rect -33361 -4420 -33301 -10
rect -33281 -4420 -33221 -10
rect -77260 -8930 -77235 -4520
rect -77215 -8930 -77155 -4520
rect -75361 -8930 -75301 -4520
rect -75281 -8930 -75256 -4520
rect -71047 -8930 -70987 -4520
rect -70967 -8930 -70907 -4520
rect -69361 -8930 -69301 -4520
rect -69281 -8930 -69221 -4520
rect -59260 -8930 -59235 -4520
rect -59215 -8930 -59155 -4520
rect -57361 -8930 -57301 -4520
rect -57281 -8930 -57221 -4520
rect -56642 -8930 -56582 -4520
rect -56562 -8930 -56502 -4520
rect -55923 -8930 -55863 -4520
rect -55843 -8930 -55783 -4520
rect -55204 -8930 -55144 -4520
rect -55124 -8930 -55064 -4520
rect -54485 -8930 -54425 -4520
rect -54405 -8930 -54345 -4520
rect -53766 -8930 -53706 -4520
rect -53686 -8930 -53626 -4520
rect -53047 -8930 -52987 -4520
rect -52967 -8930 -52907 -4520
rect -39361 -8930 -39301 -4520
rect -39281 -8930 -39221 -4520
rect -38642 -8930 -38582 -4520
rect -38562 -8930 -38502 -4520
rect -37923 -8930 -37863 -4520
rect -37843 -8930 -37783 -4520
rect -35361 -8930 -35301 -4520
rect -35281 -8930 -35221 -4520
rect -33361 -8930 -33301 -4520
rect -33281 -8930 -33221 -4520
rect -77260 -13440 -77235 -9030
rect -77215 -13440 -77155 -9030
rect -75361 -13440 -75301 -9030
rect -75281 -13440 -75256 -9030
rect -71047 -13440 -70987 -9030
rect -70967 -13440 -70907 -9030
rect -69361 -13440 -69301 -9030
rect -69281 -13440 -69221 -9030
rect -59260 -13440 -59235 -9030
rect -59215 -13440 -59155 -9030
rect -57361 -13440 -57301 -9030
rect -57281 -13440 -57221 -9030
rect -56642 -13440 -56582 -9030
rect -56562 -13440 -56502 -9030
rect -55923 -13440 -55863 -9030
rect -55843 -13440 -55783 -9030
rect -55204 -13440 -55144 -9030
rect -55124 -13440 -55064 -9030
rect -54485 -13440 -54425 -9030
rect -54405 -13440 -54345 -9030
rect -53766 -13440 -53706 -9030
rect -53686 -13440 -53626 -9030
rect -53047 -13440 -52987 -9030
rect -52967 -13440 -52907 -9030
rect -39361 -13440 -39301 -9030
rect -39281 -13440 -39221 -9030
rect -38642 -13440 -38582 -9030
rect -38562 -13440 -38502 -9030
rect -37923 -13440 -37863 -9030
rect -37843 -13440 -37783 -9030
rect -35361 -13440 -35301 -9030
rect -35281 -13440 -35221 -9030
rect -33361 -13440 -33301 -9030
rect -33281 -13440 -33221 -9030
rect -77260 -17950 -77235 -13540
rect -77215 -17950 -77155 -13540
rect -75361 -17950 -75301 -13540
rect -75281 -17950 -75256 -13540
rect -71047 -17950 -70987 -13540
rect -70967 -17950 -70907 -13540
rect -69361 -17950 -69301 -13540
rect -69281 -17950 -69221 -13540
rect -59260 -17950 -59235 -13540
rect -59215 -17950 -59155 -13540
rect -57361 -17950 -57301 -13540
rect -57281 -17950 -57221 -13540
rect -56642 -17950 -56582 -13540
rect -56562 -17950 -56502 -13540
rect -55923 -17950 -55863 -13540
rect -55843 -17950 -55783 -13540
rect -55204 -17950 -55144 -13540
rect -55124 -17950 -55064 -13540
rect -54485 -17950 -54425 -13540
rect -54405 -17950 -54345 -13540
rect -53766 -17950 -53706 -13540
rect -53686 -17950 -53626 -13540
rect -53047 -17950 -52987 -13540
rect -52967 -17950 -52907 -13540
rect -39361 -17950 -39301 -13540
rect -39281 -17950 -39221 -13540
rect -38642 -17950 -38582 -13540
rect -38562 -17950 -38502 -13540
rect -37923 -17950 -37863 -13540
rect -37843 -17950 -37783 -13540
rect -35361 -17950 -35301 -13540
rect -35281 -17950 -35221 -13540
rect -33361 -17950 -33301 -13540
rect -33281 -17950 -33221 -13540
<< error_ps >>
rect -72485 -4420 -72425 -10
rect -72405 -4420 -72345 -10
rect -71766 -4420 -71706 -10
rect -71686 -4420 -71626 -10
rect -72485 -8930 -72425 -4520
rect -72405 -8930 -72345 -4520
rect -71766 -8930 -71706 -4520
rect -71686 -8930 -71626 -4520
rect -72485 -13440 -72425 -9030
rect -72405 -13440 -72345 -9030
rect -71766 -13440 -71706 -9030
rect -71686 -13440 -71626 -9030
rect -72485 -17950 -72425 -13540
rect -72405 -17950 -72345 -13540
rect -71766 -17950 -71706 -13540
rect -71686 -17950 -71626 -13540
<< metal1 >>
rect -6400 31800 -6200 32000
rect -6400 31400 -6200 31600
rect -6400 31000 -6200 31200
rect -6400 30600 -6200 30800
rect -6400 30200 -6200 30400
rect -6400 29800 -6200 30000
rect -6400 29400 -6200 29600
rect -6400 29000 -6200 29200
rect -6400 28600 -6200 28800
rect -6400 28200 -6200 28400
rect -6400 27800 -6200 28000
rect -6400 27400 -6200 27600
rect -6400 27000 -6200 27200
rect -6400 26600 -6200 26800
rect -6400 26200 -6200 26400
rect -6400 25800 -6200 26000
rect -6400 25400 -6200 25600
rect -6400 25000 -6200 25200
rect -6400 24600 -6200 24800
rect -6400 24200 -6200 24400
rect -6400 23800 -6200 24000
rect -6400 23400 -6200 23600
rect -6400 23000 -6200 23200
rect -6400 22600 -6200 22800
rect -6400 22200 -6200 22400
rect -6400 21800 -6200 22000
rect -6400 21400 -6200 21600
rect -6400 21000 -6200 21200
rect -6400 20600 -6200 20800
rect -6400 20200 -6200 20400
rect -6400 19800 -6200 20000
rect -6400 19400 -6200 19600
rect -6400 19000 -6200 19200
rect -6400 18600 -6200 18800
rect -6400 18200 -6200 18400
rect -6400 17800 -6200 18000
rect -6400 17400 -6200 17600
rect -6400 17000 -6200 17200
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  XC1
timestamp 1665161463
transform 1 0 -64258 0 1 38040
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  XC2
timestamp 1665159686
transform 1 0 -55134 0 1 40
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  XC4
timestamp 1665159686
transform 1 0 -73134 0 1 40
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  XC5
timestamp 1665159686
transform 1 0 -38572 0 1 40
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  XC6
timestamp 1665159686
transform 1 0 -35291 0 1 38040
box -709 -18040 709 18040
use sky130_fd_pr__cap_mim_m3_1_LSQHR5  XC7
timestamp 1665159686
transform 1 0 -31650 0 1 38040
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  XC8
timestamp 1665159686
transform 1 0 -38572 0 1 38040
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  XC9
timestamp 1665159686
transform 1 0 -33291 0 1 38040
box -709 -18040 709 18040
use sky130_fd_pr__cap_mim_m3_1_EDBB5V  XC10
timestamp 1665159686
transform 1 0 -29650 0 1 38040
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_E5CB5V  XC11
timestamp 1665159686
transform 1 0 -27650 0 1 9020
box -350 -9020 349 9020
use sky130_fd_pr__cap_mim_m3_1_E9CB5V  XC12
timestamp 1665159686
transform 1 0 -21650 0 1 24510
box -350 -4510 349 4510
use sky130_fd_pr__cap_mim_m3_1_EXCB5V  XC13
timestamp 1665159686
transform 1 0 -15650 0 1 15805
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_E5CB5V  XC14
timestamp 1665159686
transform 1 0 -25650 0 1 9020
box -350 -9020 349 9020
use sky130_fd_pr__cap_mim_m3_1_E9CB5V  XC15
timestamp 1665159686
transform 1 0 -21650 0 1 13510
box -350 -4510 349 4510
use sky130_fd_pr__cap_mim_m3_1_EXCB5V  XC16
timestamp 1665159686
transform 1 0 -15650 0 1 22205
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_EXCB5V  XC17
timestamp 1665159686
transform 1 0 -17650 0 1 15805
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  XC18
timestamp 1665161463
transform 1 0 -82258 0 1 38040
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  XC19
timestamp 1665159686
transform 1 0 -55134 0 1 38040
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  XC23
timestamp 1665159686
transform 1 0 -33291 0 1 40
box -709 -18040 709 18040
use sky130_fd_pr__cap_mim_m3_1_EDBB5V  XC24
timestamp 1665159686
transform 1 0 -31650 0 1 40
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_LSQHR5  XC27
timestamp 1665159686
transform 1 0 -29650 0 1 40
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_E5CB5V  XC28
timestamp 1665159686
transform 1 0 -25650 0 1 29020
box -350 -9020 349 9020
use sky130_fd_pr__cap_mim_m3_1_E9CB5V  XC29
timestamp 1665159686
transform 1 0 -23650 0 1 13510
box -350 -4510 349 4510
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  XC30
timestamp 1665161463
transform 1 0 -17650 0 1 22205
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_E5CB5V  XC31
timestamp 1665159686
transform 1 0 -27650 0 1 29020
box -350 -9020 349 9020
use sky130_fd_pr__cap_mim_m3_1_E9CB5V  XC32
timestamp 1665159686
transform 1 0 -23650 0 1 24510
box -350 -4510 349 4510
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  XC33
timestamp 1665161463
transform 1 0 -19650 0 1 15805
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  XC34
timestamp 1665161463
transform 1 0 -19650 0 1 22205
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  sky130_fd_pr__cap_mim_m3_1_9SQ6B5_0
timestamp 1665161463
transform 1 0 -82258 0 1 40
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  sky130_fd_pr__cap_mim_m3_1_9SQ6B5_1
timestamp 1665161463
transform 1 0 -64258 0 1 40
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  sky130_fd_pr__cap_mim_m3_1_LS3JR5_0
timestamp 1665159686
transform 1 0 -42572 0 1 40
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  sky130_fd_pr__cap_mim_m3_1_LS3JR5_1
timestamp 1665159686
transform 1 0 -42572 0 1 38040
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  sky130_fd_pr__cap_mim_m3_1_LSFHR5_0
timestamp 1665159686
transform 1 0 -73134 0 1 38040
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  sky130_fd_pr__cap_mim_m3_1_LSVHR5_0
timestamp 1665159686
transform 1 0 -35291 0 1 40
box -709 -18040 709 18040
<< labels >>
flabel metal1 -6400 31800 -6200 32000 0 FreeSans 256 0 0 0 sw_sp_n9
port 0 nsew
flabel metal1 -6400 31400 -6200 31600 0 FreeSans 256 0 0 0 sw_sp_n8
port 1 nsew
flabel metal1 -6400 31000 -6200 31200 0 FreeSans 256 0 0 0 sw_sp_n7
port 2 nsew
flabel metal1 -6400 30600 -6200 30800 0 FreeSans 256 0 0 0 sw_sp_n6
port 3 nsew
flabel metal1 -6400 30200 -6200 30400 0 FreeSans 256 0 0 0 sw_sp_n5
port 4 nsew
flabel metal1 -6400 29800 -6200 30000 0 FreeSans 256 0 0 0 sw_sp_n4
port 5 nsew
flabel metal1 -6400 29400 -6200 29600 0 FreeSans 256 0 0 0 sw_sp_n3
port 6 nsew
flabel metal1 -6400 29000 -6200 29200 0 FreeSans 256 0 0 0 sw_sp_n2
port 7 nsew
flabel metal1 -6400 28600 -6200 28800 0 FreeSans 256 0 0 0 {}
port 8 nsew
flabel metal1 -6400 28200 -6200 28400 0 FreeSans 256 0 0 0 sw_sp_n1
port 9 nsew
flabel metal1 -6400 27800 -6200 28000 0 FreeSans 256 0 0 0 Vin_p
port 10 nsew
flabel metal1 -6400 27400 -6200 27600 0 FreeSans 256 0 0 0 Vin_n
port 11 nsew
flabel metal1 -6400 27000 -6200 27200 0 FreeSans 256 0 0 0 sw_sp_p9
port 12 nsew
flabel metal1 -6400 26600 -6200 26800 0 FreeSans 256 0 0 0 sw_sp_p8
port 13 nsew
flabel metal1 -6400 26200 -6200 26400 0 FreeSans 256 0 0 0 sw_sp_p7
port 14 nsew
flabel metal1 -6400 25800 -6200 26000 0 FreeSans 256 0 0 0 sw_sp_p6
port 15 nsew
flabel metal1 -6400 25400 -6200 25600 0 FreeSans 256 0 0 0 sw_sp_p5
port 16 nsew
flabel metal1 -6400 25000 -6200 25200 0 FreeSans 256 0 0 0 sw_sp_p4
port 17 nsew
flabel metal1 -6400 24600 -6200 24800 0 FreeSans 256 0 0 0 sw_sp_p3
port 18 nsew
flabel metal1 -6400 24200 -6200 24400 0 FreeSans 256 0 0 0 sw_sp_p2
port 19 nsew
flabel metal1 -6400 23800 -6200 24000 0 FreeSans 256 0 0 0 sw_sp_p1
port 20 nsew
flabel metal1 -6400 23400 -6200 23600 0 FreeSans 256 0 0 0 sw_p8
port 21 nsew
flabel metal1 -6400 23000 -6200 23200 0 FreeSans 256 0 0 0 {}
port 22 nsew
flabel metal1 -6400 22600 -6200 22800 0 FreeSans 256 0 0 0 sw_p7
port 23 nsew
flabel metal1 -6400 22200 -6200 22400 0 FreeSans 256 0 0 0 sw_p6
port 24 nsew
flabel metal1 -6400 21800 -6200 22000 0 FreeSans 256 0 0 0 sw_p5
port 25 nsew
flabel metal1 -6400 21400 -6200 21600 0 FreeSans 256 0 0 0 sw_p4
port 26 nsew
flabel metal1 -6400 21000 -6200 21200 0 FreeSans 256 0 0 0 sw_p3
port 27 nsew
flabel metal1 -6400 20600 -6200 20800 0 FreeSans 256 0 0 0 sw_p2
port 28 nsew
flabel metal1 -6400 20200 -6200 20400 0 FreeSans 256 0 0 0 sw_p1
port 29 nsew
flabel metal1 -6400 19800 -6200 20000 0 FreeSans 256 0 0 0 sw_n8
port 30 nsew
flabel metal1 -6400 19400 -6200 19600 0 FreeSans 256 0 0 0 sw_n7
port 31 nsew
flabel metal1 -6400 19000 -6200 19200 0 FreeSans 256 0 0 0 sw_n6
port 32 nsew
flabel metal1 -6400 18600 -6200 18800 0 FreeSans 256 0 0 0 sw_n5
port 33 nsew
flabel metal1 -6400 18200 -6200 18400 0 FreeSans 256 0 0 0 sw_n4
port 34 nsew
flabel metal1 -6400 17800 -6200 18000 0 FreeSans 256 0 0 0 sw_n3
port 35 nsew
flabel metal1 -6400 17400 -6200 17600 0 FreeSans 256 0 0 0 sw_n2
port 36 nsew
flabel metal1 -6400 17000 -6200 17200 0 FreeSans 256 0 0 0 sw_n1
port 37 nsew
<< end >>
