magic
tech sky130A
magscale 1 2
timestamp 1667868113
<< error_p >>
rect -791 62 -745 74
rect -599 62 -553 74
rect -407 62 -361 74
rect -215 62 -169 74
rect -23 62 23 74
rect 169 62 215 74
rect 361 62 407 74
rect 553 62 599 74
rect 745 62 791 74
rect -791 15 -785 62
rect -599 15 -593 62
rect -407 15 -401 62
rect -215 15 -209 62
rect -23 15 -17 62
rect 169 15 175 62
rect 361 15 367 62
rect 553 15 559 62
rect 745 15 751 62
rect -791 3 -745 15
rect -599 3 -553 15
rect -407 3 -361 15
rect -215 3 -169 15
rect -23 3 23 15
rect 169 3 215 15
rect 361 3 407 15
rect 553 3 599 15
rect 745 3 791 15
rect -695 -15 -649 -3
rect -503 -15 -457 -3
rect -311 -15 -265 -3
rect -119 -15 -73 -3
rect 73 -15 119 -3
rect 265 -15 311 -3
rect 457 -15 503 -3
rect 649 -15 695 -3
rect -695 -62 -689 -15
rect -503 -62 -497 -15
rect -311 -62 -305 -15
rect -119 -62 -113 -15
rect 73 -62 79 -15
rect 265 -62 271 -15
rect 457 -62 463 -15
rect 649 -62 655 -15
rect -695 -74 -649 -62
rect -503 -74 -457 -62
rect -311 -74 -265 -62
rect -119 -74 -73 -62
rect 73 -74 119 -62
rect 265 -74 311 -62
rect 457 -74 503 -62
rect 649 -74 695 -62
<< nmos >>
rect -735 -91 -705 91
rect -639 -91 -609 91
rect -543 -91 -513 91
rect -447 -91 -417 91
rect -351 -91 -321 91
rect -255 -91 -225 91
rect -159 -91 -129 91
rect -63 -91 -33 91
rect 33 -91 63 91
rect 129 -91 159 91
rect 225 -91 255 91
rect 321 -91 351 91
rect 417 -91 447 91
rect 513 -91 543 91
rect 609 -91 639 91
rect 705 -91 735 91
<< ndiff >>
rect -797 79 -735 91
rect -797 -79 -785 79
rect -751 -79 -735 79
rect -797 -91 -735 -79
rect -705 79 -639 91
rect -705 -79 -689 79
rect -655 -79 -639 79
rect -705 -91 -639 -79
rect -609 79 -543 91
rect -609 -79 -593 79
rect -559 -79 -543 79
rect -609 -91 -543 -79
rect -513 79 -447 91
rect -513 -79 -497 79
rect -463 -79 -447 79
rect -513 -91 -447 -79
rect -417 79 -351 91
rect -417 -79 -401 79
rect -367 -79 -351 79
rect -417 -91 -351 -79
rect -321 79 -255 91
rect -321 -79 -305 79
rect -271 -79 -255 79
rect -321 -91 -255 -79
rect -225 79 -159 91
rect -225 -79 -209 79
rect -175 -79 -159 79
rect -225 -91 -159 -79
rect -129 79 -63 91
rect -129 -79 -113 79
rect -79 -79 -63 79
rect -129 -91 -63 -79
rect -33 79 33 91
rect -33 -79 -17 79
rect 17 -79 33 79
rect -33 -91 33 -79
rect 63 79 129 91
rect 63 -79 79 79
rect 113 -79 129 79
rect 63 -91 129 -79
rect 159 79 225 91
rect 159 -79 175 79
rect 209 -79 225 79
rect 159 -91 225 -79
rect 255 79 321 91
rect 255 -79 271 79
rect 305 -79 321 79
rect 255 -91 321 -79
rect 351 79 417 91
rect 351 -79 367 79
rect 401 -79 417 79
rect 351 -91 417 -79
rect 447 79 513 91
rect 447 -79 463 79
rect 497 -79 513 79
rect 447 -91 513 -79
rect 543 79 609 91
rect 543 -79 559 79
rect 593 -79 609 79
rect 543 -91 609 -79
rect 639 79 705 91
rect 639 -79 655 79
rect 689 -79 705 79
rect 639 -91 705 -79
rect 735 79 797 91
rect 735 -79 751 79
rect 785 -79 797 79
rect 735 -91 797 -79
<< ndiffc >>
rect -785 -79 -751 79
rect -689 -79 -655 79
rect -593 -79 -559 79
rect -497 -79 -463 79
rect -401 -79 -367 79
rect -305 -79 -271 79
rect -209 -79 -175 79
rect -113 -79 -79 79
rect -17 -79 17 79
rect 79 -79 113 79
rect 175 -79 209 79
rect 271 -79 305 79
rect 367 -79 401 79
rect 463 -79 497 79
rect 559 -79 593 79
rect 655 -79 689 79
rect 751 -79 785 79
<< poly >>
rect -735 91 -705 121
rect -639 91 -609 121
rect -543 91 -513 121
rect -447 91 -417 121
rect -351 91 -321 121
rect -255 91 -225 121
rect -159 91 -129 121
rect -63 91 -33 121
rect 33 91 63 121
rect 129 91 159 121
rect 225 91 255 121
rect 321 91 351 121
rect 417 91 447 121
rect 513 91 543 121
rect 609 91 639 121
rect 705 91 735 121
rect -735 -113 -705 -91
rect -639 -113 -609 -91
rect -543 -113 -513 -91
rect -447 -113 -417 -91
rect -351 -113 -321 -91
rect -255 -113 -225 -91
rect -159 -113 -129 -91
rect -63 -113 -33 -91
rect 33 -113 63 -91
rect 129 -113 159 -91
rect 225 -113 255 -91
rect 321 -113 351 -91
rect 417 -113 447 -91
rect 513 -113 543 -91
rect 609 -113 639 -91
rect 705 -113 735 -91
rect -753 -129 767 -113
rect -753 -163 -737 -129
rect -703 -163 -633 -129
rect -599 -163 -545 -129
rect -511 -163 -443 -129
rect -409 -163 -353 -129
rect -319 -163 -253 -129
rect -219 -163 -161 -129
rect -127 -163 -63 -129
rect -29 -163 31 -129
rect 65 -163 127 -129
rect 161 -163 223 -129
rect 257 -163 317 -129
rect 351 -163 415 -129
rect 449 -163 507 -129
rect 541 -163 607 -129
rect 641 -163 707 -129
rect 741 -163 767 -129
rect -753 -179 767 -163
<< polycont >>
rect -737 -163 -703 -129
rect -633 -163 -599 -129
rect -545 -163 -511 -129
rect -443 -163 -409 -129
rect -353 -163 -319 -129
rect -253 -163 -219 -129
rect -161 -163 -127 -129
rect -63 -163 -29 -129
rect 31 -163 65 -129
rect 127 -163 161 -129
rect 223 -163 257 -129
rect 317 -163 351 -129
rect 415 -163 449 -129
rect 507 -163 541 -129
rect 607 -163 641 -129
rect 707 -163 741 -129
<< locali >>
rect -785 79 -751 95
rect -785 -95 -751 -79
rect -689 79 -655 95
rect -689 -95 -655 -79
rect -593 79 -559 95
rect -593 -95 -559 -79
rect -497 79 -463 95
rect -497 -95 -463 -79
rect -401 79 -367 95
rect -401 -95 -367 -79
rect -305 79 -271 95
rect -305 -95 -271 -79
rect -209 79 -175 95
rect -209 -95 -175 -79
rect -113 79 -79 95
rect -113 -95 -79 -79
rect -17 79 17 95
rect -17 -95 17 -79
rect 79 79 113 95
rect 79 -95 113 -79
rect 175 79 209 95
rect 175 -95 209 -79
rect 271 79 305 95
rect 271 -95 305 -79
rect 367 79 401 95
rect 367 -95 401 -79
rect 463 79 497 95
rect 463 -95 497 -79
rect 559 79 593 95
rect 559 -95 593 -79
rect 655 79 689 95
rect 655 -95 689 -79
rect 751 79 785 95
rect 751 -95 785 -79
rect -753 -163 -737 -129
rect -703 -163 -633 -129
rect -599 -163 -545 -129
rect -511 -163 -443 -129
rect -409 -163 -353 -129
rect -319 -163 -253 -129
rect -219 -163 -161 -129
rect -127 -163 -63 -129
rect -29 -163 31 -129
rect 65 -163 127 -129
rect 161 -163 223 -129
rect 257 -163 317 -129
rect 351 -163 415 -129
rect 449 -163 507 -129
rect 541 -163 607 -129
rect 641 -163 707 -129
rect 741 -163 767 -129
<< viali >>
rect -785 15 -751 62
rect -689 -62 -655 -15
rect -593 15 -559 62
rect -497 -62 -463 -15
rect -401 15 -367 62
rect -305 -62 -271 -15
rect -209 15 -175 62
rect -113 -62 -79 -15
rect -17 15 17 62
rect 79 -62 113 -15
rect 175 15 209 62
rect 271 -62 305 -15
rect 367 15 401 62
rect 463 -62 497 -15
rect 559 15 593 62
rect 655 -62 689 -15
rect 751 15 785 62
rect -737 -163 -703 -129
rect -633 -163 -599 -129
rect -545 -163 -511 -129
rect -443 -163 -409 -129
rect -353 -163 -319 -129
rect -253 -163 -219 -129
rect -161 -163 -127 -129
rect -63 -163 -29 -129
rect 31 -163 65 -129
rect 127 -163 161 -129
rect 223 -163 257 -129
rect 317 -163 351 -129
rect 415 -163 449 -129
rect 507 -163 541 -129
rect 607 -163 641 -129
rect 707 -163 741 -129
<< metal1 >>
rect -791 62 -745 74
rect -791 15 -785 62
rect -751 15 -745 62
rect -791 3 -745 15
rect -599 62 -553 74
rect -599 15 -593 62
rect -559 15 -553 62
rect -599 3 -553 15
rect -407 62 -361 74
rect -407 15 -401 62
rect -367 15 -361 62
rect -407 3 -361 15
rect -215 62 -169 74
rect -215 15 -209 62
rect -175 15 -169 62
rect -215 3 -169 15
rect -23 62 23 74
rect -23 15 -17 62
rect 17 15 23 62
rect -23 3 23 15
rect 169 62 215 74
rect 169 15 175 62
rect 209 15 215 62
rect 169 3 215 15
rect 361 62 407 74
rect 361 15 367 62
rect 401 15 407 62
rect 361 3 407 15
rect 553 62 599 74
rect 553 15 559 62
rect 593 15 599 62
rect 553 3 599 15
rect 745 62 791 74
rect 745 15 751 62
rect 785 15 791 62
rect 745 3 791 15
rect -695 -15 -649 -3
rect -695 -62 -689 -15
rect -655 -62 -649 -15
rect -695 -74 -649 -62
rect -503 -15 -457 -3
rect -503 -62 -497 -15
rect -463 -62 -457 -15
rect -503 -74 -457 -62
rect -311 -15 -265 -3
rect -311 -62 -305 -15
rect -271 -62 -265 -15
rect -311 -74 -265 -62
rect -119 -15 -73 -3
rect -119 -62 -113 -15
rect -79 -62 -73 -15
rect -119 -74 -73 -62
rect 73 -15 119 -3
rect 73 -62 79 -15
rect 113 -62 119 -15
rect 73 -74 119 -62
rect 265 -15 311 -3
rect 265 -62 271 -15
rect 305 -62 311 -15
rect 265 -74 311 -62
rect 457 -15 503 -3
rect 457 -62 463 -15
rect 497 -62 503 -15
rect 457 -74 503 -62
rect 649 -15 695 -3
rect 649 -62 655 -15
rect 689 -62 695 -15
rect 649 -74 695 -62
rect -753 -129 767 -123
rect -753 -163 -737 -129
rect -703 -163 -633 -129
rect -599 -163 -545 -129
rect -511 -163 -443 -129
rect -409 -163 -353 -129
rect -319 -163 -253 -129
rect -219 -163 -161 -129
rect -127 -163 -63 -129
rect -29 -163 31 -129
rect 65 -163 127 -129
rect 161 -163 223 -129
rect 257 -163 317 -129
rect 351 -163 415 -129
rect 449 -163 507 -129
rect 541 -163 607 -129
rect 641 -163 707 -129
rect 741 -163 767 -129
rect -753 -169 767 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
