magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -7976 17972 -7204 18000
rect -7976 13738 -7288 17972
rect -7224 13738 -7204 17972
rect -7976 13710 -7204 13738
rect -6964 17972 -6192 18000
rect -6964 13738 -6276 17972
rect -6212 13738 -6192 17972
rect -6964 13710 -6192 13738
rect -5952 17972 -5180 18000
rect -5952 13738 -5264 17972
rect -5200 13738 -5180 17972
rect -5952 13710 -5180 13738
rect -4940 17972 -4168 18000
rect -4940 13738 -4252 17972
rect -4188 13738 -4168 17972
rect -4940 13710 -4168 13738
rect -3928 17972 -3156 18000
rect -3928 13738 -3240 17972
rect -3176 13738 -3156 17972
rect -3928 13710 -3156 13738
rect -2916 17972 -2144 18000
rect -2916 13738 -2228 17972
rect -2164 13738 -2144 17972
rect -2916 13710 -2144 13738
rect -1904 17972 -1132 18000
rect -1904 13738 -1216 17972
rect -1152 13738 -1132 17972
rect -1904 13710 -1132 13738
rect -892 17972 -120 18000
rect -892 13738 -204 17972
rect -140 13738 -120 17972
rect -892 13710 -120 13738
rect 120 17972 892 18000
rect 120 13738 808 17972
rect 872 13738 892 17972
rect 120 13710 892 13738
rect 1132 17972 1904 18000
rect 1132 13738 1820 17972
rect 1884 13738 1904 17972
rect 1132 13710 1904 13738
rect 2144 17972 2916 18000
rect 2144 13738 2832 17972
rect 2896 13738 2916 17972
rect 2144 13710 2916 13738
rect 3156 17972 3928 18000
rect 3156 13738 3844 17972
rect 3908 13738 3928 17972
rect 3156 13710 3928 13738
rect 4168 17972 4940 18000
rect 4168 13738 4856 17972
rect 4920 13738 4940 17972
rect 4168 13710 4940 13738
rect 5180 17972 5952 18000
rect 5180 13738 5868 17972
rect 5932 13738 5952 17972
rect 5180 13710 5952 13738
rect 6192 17972 6964 18000
rect 6192 13738 6880 17972
rect 6944 13738 6964 17972
rect 6192 13710 6964 13738
rect 7204 17972 7976 18000
rect 7204 13738 7892 17972
rect 7956 13738 7976 17972
rect 7204 13710 7976 13738
rect -7976 13442 -7204 13470
rect -7976 9208 -7288 13442
rect -7224 9208 -7204 13442
rect -7976 9180 -7204 9208
rect -6964 13442 -6192 13470
rect -6964 9208 -6276 13442
rect -6212 9208 -6192 13442
rect -6964 9180 -6192 9208
rect -5952 13442 -5180 13470
rect -5952 9208 -5264 13442
rect -5200 9208 -5180 13442
rect -5952 9180 -5180 9208
rect -4940 13442 -4168 13470
rect -4940 9208 -4252 13442
rect -4188 9208 -4168 13442
rect -4940 9180 -4168 9208
rect -3928 13442 -3156 13470
rect -3928 9208 -3240 13442
rect -3176 9208 -3156 13442
rect -3928 9180 -3156 9208
rect -2916 13442 -2144 13470
rect -2916 9208 -2228 13442
rect -2164 9208 -2144 13442
rect -2916 9180 -2144 9208
rect -1904 13442 -1132 13470
rect -1904 9208 -1216 13442
rect -1152 9208 -1132 13442
rect -1904 9180 -1132 9208
rect -892 13442 -120 13470
rect -892 9208 -204 13442
rect -140 9208 -120 13442
rect -892 9180 -120 9208
rect 120 13442 892 13470
rect 120 9208 808 13442
rect 872 9208 892 13442
rect 120 9180 892 9208
rect 1132 13442 1904 13470
rect 1132 9208 1820 13442
rect 1884 9208 1904 13442
rect 1132 9180 1904 9208
rect 2144 13442 2916 13470
rect 2144 9208 2832 13442
rect 2896 9208 2916 13442
rect 2144 9180 2916 9208
rect 3156 13442 3928 13470
rect 3156 9208 3844 13442
rect 3908 9208 3928 13442
rect 3156 9180 3928 9208
rect 4168 13442 4940 13470
rect 4168 9208 4856 13442
rect 4920 9208 4940 13442
rect 4168 9180 4940 9208
rect 5180 13442 5952 13470
rect 5180 9208 5868 13442
rect 5932 9208 5952 13442
rect 5180 9180 5952 9208
rect 6192 13442 6964 13470
rect 6192 9208 6880 13442
rect 6944 9208 6964 13442
rect 6192 9180 6964 9208
rect 7204 13442 7976 13470
rect 7204 9208 7892 13442
rect 7956 9208 7976 13442
rect 7204 9180 7976 9208
rect -7976 8912 -7204 8940
rect -7976 4678 -7288 8912
rect -7224 4678 -7204 8912
rect -7976 4650 -7204 4678
rect -6964 8912 -6192 8940
rect -6964 4678 -6276 8912
rect -6212 4678 -6192 8912
rect -6964 4650 -6192 4678
rect -5952 8912 -5180 8940
rect -5952 4678 -5264 8912
rect -5200 4678 -5180 8912
rect -5952 4650 -5180 4678
rect -4940 8912 -4168 8940
rect -4940 4678 -4252 8912
rect -4188 4678 -4168 8912
rect -4940 4650 -4168 4678
rect -3928 8912 -3156 8940
rect -3928 4678 -3240 8912
rect -3176 4678 -3156 8912
rect -3928 4650 -3156 4678
rect -2916 8912 -2144 8940
rect -2916 4678 -2228 8912
rect -2164 4678 -2144 8912
rect -2916 4650 -2144 4678
rect -1904 8912 -1132 8940
rect -1904 4678 -1216 8912
rect -1152 4678 -1132 8912
rect -1904 4650 -1132 4678
rect -892 8912 -120 8940
rect -892 4678 -204 8912
rect -140 4678 -120 8912
rect -892 4650 -120 4678
rect 120 8912 892 8940
rect 120 4678 808 8912
rect 872 4678 892 8912
rect 120 4650 892 4678
rect 1132 8912 1904 8940
rect 1132 4678 1820 8912
rect 1884 4678 1904 8912
rect 1132 4650 1904 4678
rect 2144 8912 2916 8940
rect 2144 4678 2832 8912
rect 2896 4678 2916 8912
rect 2144 4650 2916 4678
rect 3156 8912 3928 8940
rect 3156 4678 3844 8912
rect 3908 4678 3928 8912
rect 3156 4650 3928 4678
rect 4168 8912 4940 8940
rect 4168 4678 4856 8912
rect 4920 4678 4940 8912
rect 4168 4650 4940 4678
rect 5180 8912 5952 8940
rect 5180 4678 5868 8912
rect 5932 4678 5952 8912
rect 5180 4650 5952 4678
rect 6192 8912 6964 8940
rect 6192 4678 6880 8912
rect 6944 4678 6964 8912
rect 6192 4650 6964 4678
rect 7204 8912 7976 8940
rect 7204 4678 7892 8912
rect 7956 4678 7976 8912
rect 7204 4650 7976 4678
rect -7976 4382 -7204 4410
rect -7976 148 -7288 4382
rect -7224 148 -7204 4382
rect -7976 120 -7204 148
rect -6964 4382 -6192 4410
rect -6964 148 -6276 4382
rect -6212 148 -6192 4382
rect -6964 120 -6192 148
rect -5952 4382 -5180 4410
rect -5952 148 -5264 4382
rect -5200 148 -5180 4382
rect -5952 120 -5180 148
rect -4940 4382 -4168 4410
rect -4940 148 -4252 4382
rect -4188 148 -4168 4382
rect -4940 120 -4168 148
rect -3928 4382 -3156 4410
rect -3928 148 -3240 4382
rect -3176 148 -3156 4382
rect -3928 120 -3156 148
rect -2916 4382 -2144 4410
rect -2916 148 -2228 4382
rect -2164 148 -2144 4382
rect -2916 120 -2144 148
rect -1904 4382 -1132 4410
rect -1904 148 -1216 4382
rect -1152 148 -1132 4382
rect -1904 120 -1132 148
rect -892 4382 -120 4410
rect -892 148 -204 4382
rect -140 148 -120 4382
rect -892 120 -120 148
rect 120 4382 892 4410
rect 120 148 808 4382
rect 872 148 892 4382
rect 120 120 892 148
rect 1132 4382 1904 4410
rect 1132 148 1820 4382
rect 1884 148 1904 4382
rect 1132 120 1904 148
rect 2144 4382 2916 4410
rect 2144 148 2832 4382
rect 2896 148 2916 4382
rect 2144 120 2916 148
rect 3156 4382 3928 4410
rect 3156 148 3844 4382
rect 3908 148 3928 4382
rect 3156 120 3928 148
rect 4168 4382 4940 4410
rect 4168 148 4856 4382
rect 4920 148 4940 4382
rect 4168 120 4940 148
rect 5180 4382 5952 4410
rect 5180 148 5868 4382
rect 5932 148 5952 4382
rect 5180 120 5952 148
rect 6192 4382 6964 4410
rect 6192 148 6880 4382
rect 6944 148 6964 4382
rect 6192 120 6964 148
rect 7204 4382 7976 4410
rect 7204 148 7892 4382
rect 7956 148 7976 4382
rect 7204 120 7976 148
rect -7976 -148 -7204 -120
rect -7976 -4382 -7288 -148
rect -7224 -4382 -7204 -148
rect -7976 -4410 -7204 -4382
rect -6964 -148 -6192 -120
rect -6964 -4382 -6276 -148
rect -6212 -4382 -6192 -148
rect -6964 -4410 -6192 -4382
rect -5952 -148 -5180 -120
rect -5952 -4382 -5264 -148
rect -5200 -4382 -5180 -148
rect -5952 -4410 -5180 -4382
rect -4940 -148 -4168 -120
rect -4940 -4382 -4252 -148
rect -4188 -4382 -4168 -148
rect -4940 -4410 -4168 -4382
rect -3928 -148 -3156 -120
rect -3928 -4382 -3240 -148
rect -3176 -4382 -3156 -148
rect -3928 -4410 -3156 -4382
rect -2916 -148 -2144 -120
rect -2916 -4382 -2228 -148
rect -2164 -4382 -2144 -148
rect -2916 -4410 -2144 -4382
rect -1904 -148 -1132 -120
rect -1904 -4382 -1216 -148
rect -1152 -4382 -1132 -148
rect -1904 -4410 -1132 -4382
rect -892 -148 -120 -120
rect -892 -4382 -204 -148
rect -140 -4382 -120 -148
rect -892 -4410 -120 -4382
rect 120 -148 892 -120
rect 120 -4382 808 -148
rect 872 -4382 892 -148
rect 120 -4410 892 -4382
rect 1132 -148 1904 -120
rect 1132 -4382 1820 -148
rect 1884 -4382 1904 -148
rect 1132 -4410 1904 -4382
rect 2144 -148 2916 -120
rect 2144 -4382 2832 -148
rect 2896 -4382 2916 -148
rect 2144 -4410 2916 -4382
rect 3156 -148 3928 -120
rect 3156 -4382 3844 -148
rect 3908 -4382 3928 -148
rect 3156 -4410 3928 -4382
rect 4168 -148 4940 -120
rect 4168 -4382 4856 -148
rect 4920 -4382 4940 -148
rect 4168 -4410 4940 -4382
rect 5180 -148 5952 -120
rect 5180 -4382 5868 -148
rect 5932 -4382 5952 -148
rect 5180 -4410 5952 -4382
rect 6192 -148 6964 -120
rect 6192 -4382 6880 -148
rect 6944 -4382 6964 -148
rect 6192 -4410 6964 -4382
rect 7204 -148 7976 -120
rect 7204 -4382 7892 -148
rect 7956 -4382 7976 -148
rect 7204 -4410 7976 -4382
rect -7976 -4678 -7204 -4650
rect -7976 -8912 -7288 -4678
rect -7224 -8912 -7204 -4678
rect -7976 -8940 -7204 -8912
rect -6964 -4678 -6192 -4650
rect -6964 -8912 -6276 -4678
rect -6212 -8912 -6192 -4678
rect -6964 -8940 -6192 -8912
rect -5952 -4678 -5180 -4650
rect -5952 -8912 -5264 -4678
rect -5200 -8912 -5180 -4678
rect -5952 -8940 -5180 -8912
rect -4940 -4678 -4168 -4650
rect -4940 -8912 -4252 -4678
rect -4188 -8912 -4168 -4678
rect -4940 -8940 -4168 -8912
rect -3928 -4678 -3156 -4650
rect -3928 -8912 -3240 -4678
rect -3176 -8912 -3156 -4678
rect -3928 -8940 -3156 -8912
rect -2916 -4678 -2144 -4650
rect -2916 -8912 -2228 -4678
rect -2164 -8912 -2144 -4678
rect -2916 -8940 -2144 -8912
rect -1904 -4678 -1132 -4650
rect -1904 -8912 -1216 -4678
rect -1152 -8912 -1132 -4678
rect -1904 -8940 -1132 -8912
rect -892 -4678 -120 -4650
rect -892 -8912 -204 -4678
rect -140 -8912 -120 -4678
rect -892 -8940 -120 -8912
rect 120 -4678 892 -4650
rect 120 -8912 808 -4678
rect 872 -8912 892 -4678
rect 120 -8940 892 -8912
rect 1132 -4678 1904 -4650
rect 1132 -8912 1820 -4678
rect 1884 -8912 1904 -4678
rect 1132 -8940 1904 -8912
rect 2144 -4678 2916 -4650
rect 2144 -8912 2832 -4678
rect 2896 -8912 2916 -4678
rect 2144 -8940 2916 -8912
rect 3156 -4678 3928 -4650
rect 3156 -8912 3844 -4678
rect 3908 -8912 3928 -4678
rect 3156 -8940 3928 -8912
rect 4168 -4678 4940 -4650
rect 4168 -8912 4856 -4678
rect 4920 -8912 4940 -4678
rect 4168 -8940 4940 -8912
rect 5180 -4678 5952 -4650
rect 5180 -8912 5868 -4678
rect 5932 -8912 5952 -4678
rect 5180 -8940 5952 -8912
rect 6192 -4678 6964 -4650
rect 6192 -8912 6880 -4678
rect 6944 -8912 6964 -4678
rect 6192 -8940 6964 -8912
rect 7204 -4678 7976 -4650
rect 7204 -8912 7892 -4678
rect 7956 -8912 7976 -4678
rect 7204 -8940 7976 -8912
rect -7976 -9208 -7204 -9180
rect -7976 -13442 -7288 -9208
rect -7224 -13442 -7204 -9208
rect -7976 -13470 -7204 -13442
rect -6964 -9208 -6192 -9180
rect -6964 -13442 -6276 -9208
rect -6212 -13442 -6192 -9208
rect -6964 -13470 -6192 -13442
rect -5952 -9208 -5180 -9180
rect -5952 -13442 -5264 -9208
rect -5200 -13442 -5180 -9208
rect -5952 -13470 -5180 -13442
rect -4940 -9208 -4168 -9180
rect -4940 -13442 -4252 -9208
rect -4188 -13442 -4168 -9208
rect -4940 -13470 -4168 -13442
rect -3928 -9208 -3156 -9180
rect -3928 -13442 -3240 -9208
rect -3176 -13442 -3156 -9208
rect -3928 -13470 -3156 -13442
rect -2916 -9208 -2144 -9180
rect -2916 -13442 -2228 -9208
rect -2164 -13442 -2144 -9208
rect -2916 -13470 -2144 -13442
rect -1904 -9208 -1132 -9180
rect -1904 -13442 -1216 -9208
rect -1152 -13442 -1132 -9208
rect -1904 -13470 -1132 -13442
rect -892 -9208 -120 -9180
rect -892 -13442 -204 -9208
rect -140 -13442 -120 -9208
rect -892 -13470 -120 -13442
rect 120 -9208 892 -9180
rect 120 -13442 808 -9208
rect 872 -13442 892 -9208
rect 120 -13470 892 -13442
rect 1132 -9208 1904 -9180
rect 1132 -13442 1820 -9208
rect 1884 -13442 1904 -9208
rect 1132 -13470 1904 -13442
rect 2144 -9208 2916 -9180
rect 2144 -13442 2832 -9208
rect 2896 -13442 2916 -9208
rect 2144 -13470 2916 -13442
rect 3156 -9208 3928 -9180
rect 3156 -13442 3844 -9208
rect 3908 -13442 3928 -9208
rect 3156 -13470 3928 -13442
rect 4168 -9208 4940 -9180
rect 4168 -13442 4856 -9208
rect 4920 -13442 4940 -9208
rect 4168 -13470 4940 -13442
rect 5180 -9208 5952 -9180
rect 5180 -13442 5868 -9208
rect 5932 -13442 5952 -9208
rect 5180 -13470 5952 -13442
rect 6192 -9208 6964 -9180
rect 6192 -13442 6880 -9208
rect 6944 -13442 6964 -9208
rect 6192 -13470 6964 -13442
rect 7204 -9208 7976 -9180
rect 7204 -13442 7892 -9208
rect 7956 -13442 7976 -9208
rect 7204 -13470 7976 -13442
rect -7976 -13738 -7204 -13710
rect -7976 -17972 -7288 -13738
rect -7224 -17972 -7204 -13738
rect -7976 -18000 -7204 -17972
rect -6964 -13738 -6192 -13710
rect -6964 -17972 -6276 -13738
rect -6212 -17972 -6192 -13738
rect -6964 -18000 -6192 -17972
rect -5952 -13738 -5180 -13710
rect -5952 -17972 -5264 -13738
rect -5200 -17972 -5180 -13738
rect -5952 -18000 -5180 -17972
rect -4940 -13738 -4168 -13710
rect -4940 -17972 -4252 -13738
rect -4188 -17972 -4168 -13738
rect -4940 -18000 -4168 -17972
rect -3928 -13738 -3156 -13710
rect -3928 -17972 -3240 -13738
rect -3176 -17972 -3156 -13738
rect -3928 -18000 -3156 -17972
rect -2916 -13738 -2144 -13710
rect -2916 -17972 -2228 -13738
rect -2164 -17972 -2144 -13738
rect -2916 -18000 -2144 -17972
rect -1904 -13738 -1132 -13710
rect -1904 -17972 -1216 -13738
rect -1152 -17972 -1132 -13738
rect -1904 -18000 -1132 -17972
rect -892 -13738 -120 -13710
rect -892 -17972 -204 -13738
rect -140 -17972 -120 -13738
rect -892 -18000 -120 -17972
rect 120 -13738 892 -13710
rect 120 -17972 808 -13738
rect 872 -17972 892 -13738
rect 120 -18000 892 -17972
rect 1132 -13738 1904 -13710
rect 1132 -17972 1820 -13738
rect 1884 -17972 1904 -13738
rect 1132 -18000 1904 -17972
rect 2144 -13738 2916 -13710
rect 2144 -17972 2832 -13738
rect 2896 -17972 2916 -13738
rect 2144 -18000 2916 -17972
rect 3156 -13738 3928 -13710
rect 3156 -17972 3844 -13738
rect 3908 -17972 3928 -13738
rect 3156 -18000 3928 -17972
rect 4168 -13738 4940 -13710
rect 4168 -17972 4856 -13738
rect 4920 -17972 4940 -13738
rect 4168 -18000 4940 -17972
rect 5180 -13738 5952 -13710
rect 5180 -17972 5868 -13738
rect 5932 -17972 5952 -13738
rect 5180 -18000 5952 -17972
rect 6192 -13738 6964 -13710
rect 6192 -17972 6880 -13738
rect 6944 -17972 6964 -13738
rect 6192 -18000 6964 -17972
rect 7204 -13738 7976 -13710
rect 7204 -17972 7892 -13738
rect 7956 -17972 7976 -13738
rect 7204 -18000 7976 -17972
<< via3 >>
rect -7288 13738 -7224 17972
rect -6276 13738 -6212 17972
rect -5264 13738 -5200 17972
rect -4252 13738 -4188 17972
rect -3240 13738 -3176 17972
rect -2228 13738 -2164 17972
rect -1216 13738 -1152 17972
rect -204 13738 -140 17972
rect 808 13738 872 17972
rect 1820 13738 1884 17972
rect 2832 13738 2896 17972
rect 3844 13738 3908 17972
rect 4856 13738 4920 17972
rect 5868 13738 5932 17972
rect 6880 13738 6944 17972
rect 7892 13738 7956 17972
rect -7288 9208 -7224 13442
rect -6276 9208 -6212 13442
rect -5264 9208 -5200 13442
rect -4252 9208 -4188 13442
rect -3240 9208 -3176 13442
rect -2228 9208 -2164 13442
rect -1216 9208 -1152 13442
rect -204 9208 -140 13442
rect 808 9208 872 13442
rect 1820 9208 1884 13442
rect 2832 9208 2896 13442
rect 3844 9208 3908 13442
rect 4856 9208 4920 13442
rect 5868 9208 5932 13442
rect 6880 9208 6944 13442
rect 7892 9208 7956 13442
rect -7288 4678 -7224 8912
rect -6276 4678 -6212 8912
rect -5264 4678 -5200 8912
rect -4252 4678 -4188 8912
rect -3240 4678 -3176 8912
rect -2228 4678 -2164 8912
rect -1216 4678 -1152 8912
rect -204 4678 -140 8912
rect 808 4678 872 8912
rect 1820 4678 1884 8912
rect 2832 4678 2896 8912
rect 3844 4678 3908 8912
rect 4856 4678 4920 8912
rect 5868 4678 5932 8912
rect 6880 4678 6944 8912
rect 7892 4678 7956 8912
rect -7288 148 -7224 4382
rect -6276 148 -6212 4382
rect -5264 148 -5200 4382
rect -4252 148 -4188 4382
rect -3240 148 -3176 4382
rect -2228 148 -2164 4382
rect -1216 148 -1152 4382
rect -204 148 -140 4382
rect 808 148 872 4382
rect 1820 148 1884 4382
rect 2832 148 2896 4382
rect 3844 148 3908 4382
rect 4856 148 4920 4382
rect 5868 148 5932 4382
rect 6880 148 6944 4382
rect 7892 148 7956 4382
rect -7288 -4382 -7224 -148
rect -6276 -4382 -6212 -148
rect -5264 -4382 -5200 -148
rect -4252 -4382 -4188 -148
rect -3240 -4382 -3176 -148
rect -2228 -4382 -2164 -148
rect -1216 -4382 -1152 -148
rect -204 -4382 -140 -148
rect 808 -4382 872 -148
rect 1820 -4382 1884 -148
rect 2832 -4382 2896 -148
rect 3844 -4382 3908 -148
rect 4856 -4382 4920 -148
rect 5868 -4382 5932 -148
rect 6880 -4382 6944 -148
rect 7892 -4382 7956 -148
rect -7288 -8912 -7224 -4678
rect -6276 -8912 -6212 -4678
rect -5264 -8912 -5200 -4678
rect -4252 -8912 -4188 -4678
rect -3240 -8912 -3176 -4678
rect -2228 -8912 -2164 -4678
rect -1216 -8912 -1152 -4678
rect -204 -8912 -140 -4678
rect 808 -8912 872 -4678
rect 1820 -8912 1884 -4678
rect 2832 -8912 2896 -4678
rect 3844 -8912 3908 -4678
rect 4856 -8912 4920 -4678
rect 5868 -8912 5932 -4678
rect 6880 -8912 6944 -4678
rect 7892 -8912 7956 -4678
rect -7288 -13442 -7224 -9208
rect -6276 -13442 -6212 -9208
rect -5264 -13442 -5200 -9208
rect -4252 -13442 -4188 -9208
rect -3240 -13442 -3176 -9208
rect -2228 -13442 -2164 -9208
rect -1216 -13442 -1152 -9208
rect -204 -13442 -140 -9208
rect 808 -13442 872 -9208
rect 1820 -13442 1884 -9208
rect 2832 -13442 2896 -9208
rect 3844 -13442 3908 -9208
rect 4856 -13442 4920 -9208
rect 5868 -13442 5932 -9208
rect 6880 -13442 6944 -9208
rect 7892 -13442 7956 -9208
rect -7288 -17972 -7224 -13738
rect -6276 -17972 -6212 -13738
rect -5264 -17972 -5200 -13738
rect -4252 -17972 -4188 -13738
rect -3240 -17972 -3176 -13738
rect -2228 -17972 -2164 -13738
rect -1216 -17972 -1152 -13738
rect -204 -17972 -140 -13738
rect 808 -17972 872 -13738
rect 1820 -17972 1884 -13738
rect 2832 -17972 2896 -13738
rect 3844 -17972 3908 -13738
rect 4856 -17972 4920 -13738
rect 5868 -17972 5932 -13738
rect 6880 -17972 6944 -13738
rect 7892 -17972 7956 -13738
<< mimcap >>
rect -7936 17920 -7536 17960
rect -7936 13790 -7896 17920
rect -7576 13790 -7536 17920
rect -7936 13750 -7536 13790
rect -6924 17920 -6524 17960
rect -6924 13790 -6884 17920
rect -6564 13790 -6524 17920
rect -6924 13750 -6524 13790
rect -5912 17920 -5512 17960
rect -5912 13790 -5872 17920
rect -5552 13790 -5512 17920
rect -5912 13750 -5512 13790
rect -4900 17920 -4500 17960
rect -4900 13790 -4860 17920
rect -4540 13790 -4500 17920
rect -4900 13750 -4500 13790
rect -3888 17920 -3488 17960
rect -3888 13790 -3848 17920
rect -3528 13790 -3488 17920
rect -3888 13750 -3488 13790
rect -2876 17920 -2476 17960
rect -2876 13790 -2836 17920
rect -2516 13790 -2476 17920
rect -2876 13750 -2476 13790
rect -1864 17920 -1464 17960
rect -1864 13790 -1824 17920
rect -1504 13790 -1464 17920
rect -1864 13750 -1464 13790
rect -852 17920 -452 17960
rect -852 13790 -812 17920
rect -492 13790 -452 17920
rect -852 13750 -452 13790
rect 160 17920 560 17960
rect 160 13790 200 17920
rect 520 13790 560 17920
rect 160 13750 560 13790
rect 1172 17920 1572 17960
rect 1172 13790 1212 17920
rect 1532 13790 1572 17920
rect 1172 13750 1572 13790
rect 2184 17920 2584 17960
rect 2184 13790 2224 17920
rect 2544 13790 2584 17920
rect 2184 13750 2584 13790
rect 3196 17920 3596 17960
rect 3196 13790 3236 17920
rect 3556 13790 3596 17920
rect 3196 13750 3596 13790
rect 4208 17920 4608 17960
rect 4208 13790 4248 17920
rect 4568 13790 4608 17920
rect 4208 13750 4608 13790
rect 5220 17920 5620 17960
rect 5220 13790 5260 17920
rect 5580 13790 5620 17920
rect 5220 13750 5620 13790
rect 6232 17920 6632 17960
rect 6232 13790 6272 17920
rect 6592 13790 6632 17920
rect 6232 13750 6632 13790
rect 7244 17920 7644 17960
rect 7244 13790 7284 17920
rect 7604 13790 7644 17920
rect 7244 13750 7644 13790
rect -7936 13390 -7536 13430
rect -7936 9260 -7896 13390
rect -7576 9260 -7536 13390
rect -7936 9220 -7536 9260
rect -6924 13390 -6524 13430
rect -6924 9260 -6884 13390
rect -6564 9260 -6524 13390
rect -6924 9220 -6524 9260
rect -5912 13390 -5512 13430
rect -5912 9260 -5872 13390
rect -5552 9260 -5512 13390
rect -5912 9220 -5512 9260
rect -4900 13390 -4500 13430
rect -4900 9260 -4860 13390
rect -4540 9260 -4500 13390
rect -4900 9220 -4500 9260
rect -3888 13390 -3488 13430
rect -3888 9260 -3848 13390
rect -3528 9260 -3488 13390
rect -3888 9220 -3488 9260
rect -2876 13390 -2476 13430
rect -2876 9260 -2836 13390
rect -2516 9260 -2476 13390
rect -2876 9220 -2476 9260
rect -1864 13390 -1464 13430
rect -1864 9260 -1824 13390
rect -1504 9260 -1464 13390
rect -1864 9220 -1464 9260
rect -852 13390 -452 13430
rect -852 9260 -812 13390
rect -492 9260 -452 13390
rect -852 9220 -452 9260
rect 160 13390 560 13430
rect 160 9260 200 13390
rect 520 9260 560 13390
rect 160 9220 560 9260
rect 1172 13390 1572 13430
rect 1172 9260 1212 13390
rect 1532 9260 1572 13390
rect 1172 9220 1572 9260
rect 2184 13390 2584 13430
rect 2184 9260 2224 13390
rect 2544 9260 2584 13390
rect 2184 9220 2584 9260
rect 3196 13390 3596 13430
rect 3196 9260 3236 13390
rect 3556 9260 3596 13390
rect 3196 9220 3596 9260
rect 4208 13390 4608 13430
rect 4208 9260 4248 13390
rect 4568 9260 4608 13390
rect 4208 9220 4608 9260
rect 5220 13390 5620 13430
rect 5220 9260 5260 13390
rect 5580 9260 5620 13390
rect 5220 9220 5620 9260
rect 6232 13390 6632 13430
rect 6232 9260 6272 13390
rect 6592 9260 6632 13390
rect 6232 9220 6632 9260
rect 7244 13390 7644 13430
rect 7244 9260 7284 13390
rect 7604 9260 7644 13390
rect 7244 9220 7644 9260
rect -7936 8860 -7536 8900
rect -7936 4730 -7896 8860
rect -7576 4730 -7536 8860
rect -7936 4690 -7536 4730
rect -6924 8860 -6524 8900
rect -6924 4730 -6884 8860
rect -6564 4730 -6524 8860
rect -6924 4690 -6524 4730
rect -5912 8860 -5512 8900
rect -5912 4730 -5872 8860
rect -5552 4730 -5512 8860
rect -5912 4690 -5512 4730
rect -4900 8860 -4500 8900
rect -4900 4730 -4860 8860
rect -4540 4730 -4500 8860
rect -4900 4690 -4500 4730
rect -3888 8860 -3488 8900
rect -3888 4730 -3848 8860
rect -3528 4730 -3488 8860
rect -3888 4690 -3488 4730
rect -2876 8860 -2476 8900
rect -2876 4730 -2836 8860
rect -2516 4730 -2476 8860
rect -2876 4690 -2476 4730
rect -1864 8860 -1464 8900
rect -1864 4730 -1824 8860
rect -1504 4730 -1464 8860
rect -1864 4690 -1464 4730
rect -852 8860 -452 8900
rect -852 4730 -812 8860
rect -492 4730 -452 8860
rect -852 4690 -452 4730
rect 160 8860 560 8900
rect 160 4730 200 8860
rect 520 4730 560 8860
rect 160 4690 560 4730
rect 1172 8860 1572 8900
rect 1172 4730 1212 8860
rect 1532 4730 1572 8860
rect 1172 4690 1572 4730
rect 2184 8860 2584 8900
rect 2184 4730 2224 8860
rect 2544 4730 2584 8860
rect 2184 4690 2584 4730
rect 3196 8860 3596 8900
rect 3196 4730 3236 8860
rect 3556 4730 3596 8860
rect 3196 4690 3596 4730
rect 4208 8860 4608 8900
rect 4208 4730 4248 8860
rect 4568 4730 4608 8860
rect 4208 4690 4608 4730
rect 5220 8860 5620 8900
rect 5220 4730 5260 8860
rect 5580 4730 5620 8860
rect 5220 4690 5620 4730
rect 6232 8860 6632 8900
rect 6232 4730 6272 8860
rect 6592 4730 6632 8860
rect 6232 4690 6632 4730
rect 7244 8860 7644 8900
rect 7244 4730 7284 8860
rect 7604 4730 7644 8860
rect 7244 4690 7644 4730
rect -7936 4330 -7536 4370
rect -7936 200 -7896 4330
rect -7576 200 -7536 4330
rect -7936 160 -7536 200
rect -6924 4330 -6524 4370
rect -6924 200 -6884 4330
rect -6564 200 -6524 4330
rect -6924 160 -6524 200
rect -5912 4330 -5512 4370
rect -5912 200 -5872 4330
rect -5552 200 -5512 4330
rect -5912 160 -5512 200
rect -4900 4330 -4500 4370
rect -4900 200 -4860 4330
rect -4540 200 -4500 4330
rect -4900 160 -4500 200
rect -3888 4330 -3488 4370
rect -3888 200 -3848 4330
rect -3528 200 -3488 4330
rect -3888 160 -3488 200
rect -2876 4330 -2476 4370
rect -2876 200 -2836 4330
rect -2516 200 -2476 4330
rect -2876 160 -2476 200
rect -1864 4330 -1464 4370
rect -1864 200 -1824 4330
rect -1504 200 -1464 4330
rect -1864 160 -1464 200
rect -852 4330 -452 4370
rect -852 200 -812 4330
rect -492 200 -452 4330
rect -852 160 -452 200
rect 160 4330 560 4370
rect 160 200 200 4330
rect 520 200 560 4330
rect 160 160 560 200
rect 1172 4330 1572 4370
rect 1172 200 1212 4330
rect 1532 200 1572 4330
rect 1172 160 1572 200
rect 2184 4330 2584 4370
rect 2184 200 2224 4330
rect 2544 200 2584 4330
rect 2184 160 2584 200
rect 3196 4330 3596 4370
rect 3196 200 3236 4330
rect 3556 200 3596 4330
rect 3196 160 3596 200
rect 4208 4330 4608 4370
rect 4208 200 4248 4330
rect 4568 200 4608 4330
rect 4208 160 4608 200
rect 5220 4330 5620 4370
rect 5220 200 5260 4330
rect 5580 200 5620 4330
rect 5220 160 5620 200
rect 6232 4330 6632 4370
rect 6232 200 6272 4330
rect 6592 200 6632 4330
rect 6232 160 6632 200
rect 7244 4330 7644 4370
rect 7244 200 7284 4330
rect 7604 200 7644 4330
rect 7244 160 7644 200
rect -7936 -200 -7536 -160
rect -7936 -4330 -7896 -200
rect -7576 -4330 -7536 -200
rect -7936 -4370 -7536 -4330
rect -6924 -200 -6524 -160
rect -6924 -4330 -6884 -200
rect -6564 -4330 -6524 -200
rect -6924 -4370 -6524 -4330
rect -5912 -200 -5512 -160
rect -5912 -4330 -5872 -200
rect -5552 -4330 -5512 -200
rect -5912 -4370 -5512 -4330
rect -4900 -200 -4500 -160
rect -4900 -4330 -4860 -200
rect -4540 -4330 -4500 -200
rect -4900 -4370 -4500 -4330
rect -3888 -200 -3488 -160
rect -3888 -4330 -3848 -200
rect -3528 -4330 -3488 -200
rect -3888 -4370 -3488 -4330
rect -2876 -200 -2476 -160
rect -2876 -4330 -2836 -200
rect -2516 -4330 -2476 -200
rect -2876 -4370 -2476 -4330
rect -1864 -200 -1464 -160
rect -1864 -4330 -1824 -200
rect -1504 -4330 -1464 -200
rect -1864 -4370 -1464 -4330
rect -852 -200 -452 -160
rect -852 -4330 -812 -200
rect -492 -4330 -452 -200
rect -852 -4370 -452 -4330
rect 160 -200 560 -160
rect 160 -4330 200 -200
rect 520 -4330 560 -200
rect 160 -4370 560 -4330
rect 1172 -200 1572 -160
rect 1172 -4330 1212 -200
rect 1532 -4330 1572 -200
rect 1172 -4370 1572 -4330
rect 2184 -200 2584 -160
rect 2184 -4330 2224 -200
rect 2544 -4330 2584 -200
rect 2184 -4370 2584 -4330
rect 3196 -200 3596 -160
rect 3196 -4330 3236 -200
rect 3556 -4330 3596 -200
rect 3196 -4370 3596 -4330
rect 4208 -200 4608 -160
rect 4208 -4330 4248 -200
rect 4568 -4330 4608 -200
rect 4208 -4370 4608 -4330
rect 5220 -200 5620 -160
rect 5220 -4330 5260 -200
rect 5580 -4330 5620 -200
rect 5220 -4370 5620 -4330
rect 6232 -200 6632 -160
rect 6232 -4330 6272 -200
rect 6592 -4330 6632 -200
rect 6232 -4370 6632 -4330
rect 7244 -200 7644 -160
rect 7244 -4330 7284 -200
rect 7604 -4330 7644 -200
rect 7244 -4370 7644 -4330
rect -7936 -4730 -7536 -4690
rect -7936 -8860 -7896 -4730
rect -7576 -8860 -7536 -4730
rect -7936 -8900 -7536 -8860
rect -6924 -4730 -6524 -4690
rect -6924 -8860 -6884 -4730
rect -6564 -8860 -6524 -4730
rect -6924 -8900 -6524 -8860
rect -5912 -4730 -5512 -4690
rect -5912 -8860 -5872 -4730
rect -5552 -8860 -5512 -4730
rect -5912 -8900 -5512 -8860
rect -4900 -4730 -4500 -4690
rect -4900 -8860 -4860 -4730
rect -4540 -8860 -4500 -4730
rect -4900 -8900 -4500 -8860
rect -3888 -4730 -3488 -4690
rect -3888 -8860 -3848 -4730
rect -3528 -8860 -3488 -4730
rect -3888 -8900 -3488 -8860
rect -2876 -4730 -2476 -4690
rect -2876 -8860 -2836 -4730
rect -2516 -8860 -2476 -4730
rect -2876 -8900 -2476 -8860
rect -1864 -4730 -1464 -4690
rect -1864 -8860 -1824 -4730
rect -1504 -8860 -1464 -4730
rect -1864 -8900 -1464 -8860
rect -852 -4730 -452 -4690
rect -852 -8860 -812 -4730
rect -492 -8860 -452 -4730
rect -852 -8900 -452 -8860
rect 160 -4730 560 -4690
rect 160 -8860 200 -4730
rect 520 -8860 560 -4730
rect 160 -8900 560 -8860
rect 1172 -4730 1572 -4690
rect 1172 -8860 1212 -4730
rect 1532 -8860 1572 -4730
rect 1172 -8900 1572 -8860
rect 2184 -4730 2584 -4690
rect 2184 -8860 2224 -4730
rect 2544 -8860 2584 -4730
rect 2184 -8900 2584 -8860
rect 3196 -4730 3596 -4690
rect 3196 -8860 3236 -4730
rect 3556 -8860 3596 -4730
rect 3196 -8900 3596 -8860
rect 4208 -4730 4608 -4690
rect 4208 -8860 4248 -4730
rect 4568 -8860 4608 -4730
rect 4208 -8900 4608 -8860
rect 5220 -4730 5620 -4690
rect 5220 -8860 5260 -4730
rect 5580 -8860 5620 -4730
rect 5220 -8900 5620 -8860
rect 6232 -4730 6632 -4690
rect 6232 -8860 6272 -4730
rect 6592 -8860 6632 -4730
rect 6232 -8900 6632 -8860
rect 7244 -4730 7644 -4690
rect 7244 -8860 7284 -4730
rect 7604 -8860 7644 -4730
rect 7244 -8900 7644 -8860
rect -7936 -9260 -7536 -9220
rect -7936 -13390 -7896 -9260
rect -7576 -13390 -7536 -9260
rect -7936 -13430 -7536 -13390
rect -6924 -9260 -6524 -9220
rect -6924 -13390 -6884 -9260
rect -6564 -13390 -6524 -9260
rect -6924 -13430 -6524 -13390
rect -5912 -9260 -5512 -9220
rect -5912 -13390 -5872 -9260
rect -5552 -13390 -5512 -9260
rect -5912 -13430 -5512 -13390
rect -4900 -9260 -4500 -9220
rect -4900 -13390 -4860 -9260
rect -4540 -13390 -4500 -9260
rect -4900 -13430 -4500 -13390
rect -3888 -9260 -3488 -9220
rect -3888 -13390 -3848 -9260
rect -3528 -13390 -3488 -9260
rect -3888 -13430 -3488 -13390
rect -2876 -9260 -2476 -9220
rect -2876 -13390 -2836 -9260
rect -2516 -13390 -2476 -9260
rect -2876 -13430 -2476 -13390
rect -1864 -9260 -1464 -9220
rect -1864 -13390 -1824 -9260
rect -1504 -13390 -1464 -9260
rect -1864 -13430 -1464 -13390
rect -852 -9260 -452 -9220
rect -852 -13390 -812 -9260
rect -492 -13390 -452 -9260
rect -852 -13430 -452 -13390
rect 160 -9260 560 -9220
rect 160 -13390 200 -9260
rect 520 -13390 560 -9260
rect 160 -13430 560 -13390
rect 1172 -9260 1572 -9220
rect 1172 -13390 1212 -9260
rect 1532 -13390 1572 -9260
rect 1172 -13430 1572 -13390
rect 2184 -9260 2584 -9220
rect 2184 -13390 2224 -9260
rect 2544 -13390 2584 -9260
rect 2184 -13430 2584 -13390
rect 3196 -9260 3596 -9220
rect 3196 -13390 3236 -9260
rect 3556 -13390 3596 -9260
rect 3196 -13430 3596 -13390
rect 4208 -9260 4608 -9220
rect 4208 -13390 4248 -9260
rect 4568 -13390 4608 -9260
rect 4208 -13430 4608 -13390
rect 5220 -9260 5620 -9220
rect 5220 -13390 5260 -9260
rect 5580 -13390 5620 -9260
rect 5220 -13430 5620 -13390
rect 6232 -9260 6632 -9220
rect 6232 -13390 6272 -9260
rect 6592 -13390 6632 -9260
rect 6232 -13430 6632 -13390
rect 7244 -9260 7644 -9220
rect 7244 -13390 7284 -9260
rect 7604 -13390 7644 -9260
rect 7244 -13430 7644 -13390
rect -7936 -13790 -7536 -13750
rect -7936 -17920 -7896 -13790
rect -7576 -17920 -7536 -13790
rect -7936 -17960 -7536 -17920
rect -6924 -13790 -6524 -13750
rect -6924 -17920 -6884 -13790
rect -6564 -17920 -6524 -13790
rect -6924 -17960 -6524 -17920
rect -5912 -13790 -5512 -13750
rect -5912 -17920 -5872 -13790
rect -5552 -17920 -5512 -13790
rect -5912 -17960 -5512 -17920
rect -4900 -13790 -4500 -13750
rect -4900 -17920 -4860 -13790
rect -4540 -17920 -4500 -13790
rect -4900 -17960 -4500 -17920
rect -3888 -13790 -3488 -13750
rect -3888 -17920 -3848 -13790
rect -3528 -17920 -3488 -13790
rect -3888 -17960 -3488 -17920
rect -2876 -13790 -2476 -13750
rect -2876 -17920 -2836 -13790
rect -2516 -17920 -2476 -13790
rect -2876 -17960 -2476 -17920
rect -1864 -13790 -1464 -13750
rect -1864 -17920 -1824 -13790
rect -1504 -17920 -1464 -13790
rect -1864 -17960 -1464 -17920
rect -852 -13790 -452 -13750
rect -852 -17920 -812 -13790
rect -492 -17920 -452 -13790
rect -852 -17960 -452 -17920
rect 160 -13790 560 -13750
rect 160 -17920 200 -13790
rect 520 -17920 560 -13790
rect 160 -17960 560 -17920
rect 1172 -13790 1572 -13750
rect 1172 -17920 1212 -13790
rect 1532 -17920 1572 -13790
rect 1172 -17960 1572 -17920
rect 2184 -13790 2584 -13750
rect 2184 -17920 2224 -13790
rect 2544 -17920 2584 -13790
rect 2184 -17960 2584 -17920
rect 3196 -13790 3596 -13750
rect 3196 -17920 3236 -13790
rect 3556 -17920 3596 -13790
rect 3196 -17960 3596 -17920
rect 4208 -13790 4608 -13750
rect 4208 -17920 4248 -13790
rect 4568 -17920 4608 -13790
rect 4208 -17960 4608 -17920
rect 5220 -13790 5620 -13750
rect 5220 -17920 5260 -13790
rect 5580 -17920 5620 -13790
rect 5220 -17960 5620 -17920
rect 6232 -13790 6632 -13750
rect 6232 -17920 6272 -13790
rect 6592 -17920 6632 -13790
rect 6232 -17960 6632 -17920
rect 7244 -13790 7644 -13750
rect 7244 -17920 7284 -13790
rect 7604 -17920 7644 -13790
rect 7244 -17960 7644 -17920
<< mimcapcontact >>
rect -7896 13790 -7576 17920
rect -6884 13790 -6564 17920
rect -5872 13790 -5552 17920
rect -4860 13790 -4540 17920
rect -3848 13790 -3528 17920
rect -2836 13790 -2516 17920
rect -1824 13790 -1504 17920
rect -812 13790 -492 17920
rect 200 13790 520 17920
rect 1212 13790 1532 17920
rect 2224 13790 2544 17920
rect 3236 13790 3556 17920
rect 4248 13790 4568 17920
rect 5260 13790 5580 17920
rect 6272 13790 6592 17920
rect 7284 13790 7604 17920
rect -7896 9260 -7576 13390
rect -6884 9260 -6564 13390
rect -5872 9260 -5552 13390
rect -4860 9260 -4540 13390
rect -3848 9260 -3528 13390
rect -2836 9260 -2516 13390
rect -1824 9260 -1504 13390
rect -812 9260 -492 13390
rect 200 9260 520 13390
rect 1212 9260 1532 13390
rect 2224 9260 2544 13390
rect 3236 9260 3556 13390
rect 4248 9260 4568 13390
rect 5260 9260 5580 13390
rect 6272 9260 6592 13390
rect 7284 9260 7604 13390
rect -7896 4730 -7576 8860
rect -6884 4730 -6564 8860
rect -5872 4730 -5552 8860
rect -4860 4730 -4540 8860
rect -3848 4730 -3528 8860
rect -2836 4730 -2516 8860
rect -1824 4730 -1504 8860
rect -812 4730 -492 8860
rect 200 4730 520 8860
rect 1212 4730 1532 8860
rect 2224 4730 2544 8860
rect 3236 4730 3556 8860
rect 4248 4730 4568 8860
rect 5260 4730 5580 8860
rect 6272 4730 6592 8860
rect 7284 4730 7604 8860
rect -7896 200 -7576 4330
rect -6884 200 -6564 4330
rect -5872 200 -5552 4330
rect -4860 200 -4540 4330
rect -3848 200 -3528 4330
rect -2836 200 -2516 4330
rect -1824 200 -1504 4330
rect -812 200 -492 4330
rect 200 200 520 4330
rect 1212 200 1532 4330
rect 2224 200 2544 4330
rect 3236 200 3556 4330
rect 4248 200 4568 4330
rect 5260 200 5580 4330
rect 6272 200 6592 4330
rect 7284 200 7604 4330
rect -7896 -4330 -7576 -200
rect -6884 -4330 -6564 -200
rect -5872 -4330 -5552 -200
rect -4860 -4330 -4540 -200
rect -3848 -4330 -3528 -200
rect -2836 -4330 -2516 -200
rect -1824 -4330 -1504 -200
rect -812 -4330 -492 -200
rect 200 -4330 520 -200
rect 1212 -4330 1532 -200
rect 2224 -4330 2544 -200
rect 3236 -4330 3556 -200
rect 4248 -4330 4568 -200
rect 5260 -4330 5580 -200
rect 6272 -4330 6592 -200
rect 7284 -4330 7604 -200
rect -7896 -8860 -7576 -4730
rect -6884 -8860 -6564 -4730
rect -5872 -8860 -5552 -4730
rect -4860 -8860 -4540 -4730
rect -3848 -8860 -3528 -4730
rect -2836 -8860 -2516 -4730
rect -1824 -8860 -1504 -4730
rect -812 -8860 -492 -4730
rect 200 -8860 520 -4730
rect 1212 -8860 1532 -4730
rect 2224 -8860 2544 -4730
rect 3236 -8860 3556 -4730
rect 4248 -8860 4568 -4730
rect 5260 -8860 5580 -4730
rect 6272 -8860 6592 -4730
rect 7284 -8860 7604 -4730
rect -7896 -13390 -7576 -9260
rect -6884 -13390 -6564 -9260
rect -5872 -13390 -5552 -9260
rect -4860 -13390 -4540 -9260
rect -3848 -13390 -3528 -9260
rect -2836 -13390 -2516 -9260
rect -1824 -13390 -1504 -9260
rect -812 -13390 -492 -9260
rect 200 -13390 520 -9260
rect 1212 -13390 1532 -9260
rect 2224 -13390 2544 -9260
rect 3236 -13390 3556 -9260
rect 4248 -13390 4568 -9260
rect 5260 -13390 5580 -9260
rect 6272 -13390 6592 -9260
rect 7284 -13390 7604 -9260
rect -7896 -17920 -7576 -13790
rect -6884 -17920 -6564 -13790
rect -5872 -17920 -5552 -13790
rect -4860 -17920 -4540 -13790
rect -3848 -17920 -3528 -13790
rect -2836 -17920 -2516 -13790
rect -1824 -17920 -1504 -13790
rect -812 -17920 -492 -13790
rect 200 -17920 520 -13790
rect 1212 -17920 1532 -13790
rect 2224 -17920 2544 -13790
rect 3236 -17920 3556 -13790
rect 4248 -17920 4568 -13790
rect 5260 -17920 5580 -13790
rect 6272 -17920 6592 -13790
rect 7284 -17920 7604 -13790
<< metal4 >>
rect -7788 17921 -7684 18120
rect -7308 17972 -7204 18120
rect -7897 17920 -7575 17921
rect -7897 13790 -7896 17920
rect -7576 13790 -7575 17920
rect -7897 13789 -7575 13790
rect -7788 13391 -7684 13789
rect -7308 13738 -7288 17972
rect -7224 13738 -7204 17972
rect -6776 17921 -6672 18120
rect -6296 17972 -6192 18120
rect -6885 17920 -6563 17921
rect -6885 13790 -6884 17920
rect -6564 13790 -6563 17920
rect -6885 13789 -6563 13790
rect -7308 13442 -7204 13738
rect -7897 13390 -7575 13391
rect -7897 9260 -7896 13390
rect -7576 9260 -7575 13390
rect -7897 9259 -7575 9260
rect -7788 8861 -7684 9259
rect -7308 9208 -7288 13442
rect -7224 9208 -7204 13442
rect -6776 13391 -6672 13789
rect -6296 13738 -6276 17972
rect -6212 13738 -6192 17972
rect -5764 17921 -5660 18120
rect -5284 17972 -5180 18120
rect -5873 17920 -5551 17921
rect -5873 13790 -5872 17920
rect -5552 13790 -5551 17920
rect -5873 13789 -5551 13790
rect -6296 13442 -6192 13738
rect -6885 13390 -6563 13391
rect -6885 9260 -6884 13390
rect -6564 9260 -6563 13390
rect -6885 9259 -6563 9260
rect -7308 8912 -7204 9208
rect -7897 8860 -7575 8861
rect -7897 4730 -7896 8860
rect -7576 4730 -7575 8860
rect -7897 4729 -7575 4730
rect -7788 4331 -7684 4729
rect -7308 4678 -7288 8912
rect -7224 4678 -7204 8912
rect -6776 8861 -6672 9259
rect -6296 9208 -6276 13442
rect -6212 9208 -6192 13442
rect -5764 13391 -5660 13789
rect -5284 13738 -5264 17972
rect -5200 13738 -5180 17972
rect -4752 17921 -4648 18120
rect -4272 17972 -4168 18120
rect -4861 17920 -4539 17921
rect -4861 13790 -4860 17920
rect -4540 13790 -4539 17920
rect -4861 13789 -4539 13790
rect -5284 13442 -5180 13738
rect -5873 13390 -5551 13391
rect -5873 9260 -5872 13390
rect -5552 9260 -5551 13390
rect -5873 9259 -5551 9260
rect -6296 8912 -6192 9208
rect -6885 8860 -6563 8861
rect -6885 4730 -6884 8860
rect -6564 4730 -6563 8860
rect -6885 4729 -6563 4730
rect -7308 4382 -7204 4678
rect -7897 4330 -7575 4331
rect -7897 200 -7896 4330
rect -7576 200 -7575 4330
rect -7897 199 -7575 200
rect -7788 -199 -7684 199
rect -7308 148 -7288 4382
rect -7224 148 -7204 4382
rect -6776 4331 -6672 4729
rect -6296 4678 -6276 8912
rect -6212 4678 -6192 8912
rect -5764 8861 -5660 9259
rect -5284 9208 -5264 13442
rect -5200 9208 -5180 13442
rect -4752 13391 -4648 13789
rect -4272 13738 -4252 17972
rect -4188 13738 -4168 17972
rect -3740 17921 -3636 18120
rect -3260 17972 -3156 18120
rect -3849 17920 -3527 17921
rect -3849 13790 -3848 17920
rect -3528 13790 -3527 17920
rect -3849 13789 -3527 13790
rect -4272 13442 -4168 13738
rect -4861 13390 -4539 13391
rect -4861 9260 -4860 13390
rect -4540 9260 -4539 13390
rect -4861 9259 -4539 9260
rect -5284 8912 -5180 9208
rect -5873 8860 -5551 8861
rect -5873 4730 -5872 8860
rect -5552 4730 -5551 8860
rect -5873 4729 -5551 4730
rect -6296 4382 -6192 4678
rect -6885 4330 -6563 4331
rect -6885 200 -6884 4330
rect -6564 200 -6563 4330
rect -6885 199 -6563 200
rect -7308 -148 -7204 148
rect -7897 -200 -7575 -199
rect -7897 -4330 -7896 -200
rect -7576 -4330 -7575 -200
rect -7897 -4331 -7575 -4330
rect -7788 -4729 -7684 -4331
rect -7308 -4382 -7288 -148
rect -7224 -4382 -7204 -148
rect -6776 -199 -6672 199
rect -6296 148 -6276 4382
rect -6212 148 -6192 4382
rect -5764 4331 -5660 4729
rect -5284 4678 -5264 8912
rect -5200 4678 -5180 8912
rect -4752 8861 -4648 9259
rect -4272 9208 -4252 13442
rect -4188 9208 -4168 13442
rect -3740 13391 -3636 13789
rect -3260 13738 -3240 17972
rect -3176 13738 -3156 17972
rect -2728 17921 -2624 18120
rect -2248 17972 -2144 18120
rect -2837 17920 -2515 17921
rect -2837 13790 -2836 17920
rect -2516 13790 -2515 17920
rect -2837 13789 -2515 13790
rect -3260 13442 -3156 13738
rect -3849 13390 -3527 13391
rect -3849 9260 -3848 13390
rect -3528 9260 -3527 13390
rect -3849 9259 -3527 9260
rect -4272 8912 -4168 9208
rect -4861 8860 -4539 8861
rect -4861 4730 -4860 8860
rect -4540 4730 -4539 8860
rect -4861 4729 -4539 4730
rect -5284 4382 -5180 4678
rect -5873 4330 -5551 4331
rect -5873 200 -5872 4330
rect -5552 200 -5551 4330
rect -5873 199 -5551 200
rect -6296 -148 -6192 148
rect -6885 -200 -6563 -199
rect -6885 -4330 -6884 -200
rect -6564 -4330 -6563 -200
rect -6885 -4331 -6563 -4330
rect -7308 -4678 -7204 -4382
rect -7897 -4730 -7575 -4729
rect -7897 -8860 -7896 -4730
rect -7576 -8860 -7575 -4730
rect -7897 -8861 -7575 -8860
rect -7788 -9259 -7684 -8861
rect -7308 -8912 -7288 -4678
rect -7224 -8912 -7204 -4678
rect -6776 -4729 -6672 -4331
rect -6296 -4382 -6276 -148
rect -6212 -4382 -6192 -148
rect -5764 -199 -5660 199
rect -5284 148 -5264 4382
rect -5200 148 -5180 4382
rect -4752 4331 -4648 4729
rect -4272 4678 -4252 8912
rect -4188 4678 -4168 8912
rect -3740 8861 -3636 9259
rect -3260 9208 -3240 13442
rect -3176 9208 -3156 13442
rect -2728 13391 -2624 13789
rect -2248 13738 -2228 17972
rect -2164 13738 -2144 17972
rect -1716 17921 -1612 18120
rect -1236 17972 -1132 18120
rect -1825 17920 -1503 17921
rect -1825 13790 -1824 17920
rect -1504 13790 -1503 17920
rect -1825 13789 -1503 13790
rect -2248 13442 -2144 13738
rect -2837 13390 -2515 13391
rect -2837 9260 -2836 13390
rect -2516 9260 -2515 13390
rect -2837 9259 -2515 9260
rect -3260 8912 -3156 9208
rect -3849 8860 -3527 8861
rect -3849 4730 -3848 8860
rect -3528 4730 -3527 8860
rect -3849 4729 -3527 4730
rect -4272 4382 -4168 4678
rect -4861 4330 -4539 4331
rect -4861 200 -4860 4330
rect -4540 200 -4539 4330
rect -4861 199 -4539 200
rect -5284 -148 -5180 148
rect -5873 -200 -5551 -199
rect -5873 -4330 -5872 -200
rect -5552 -4330 -5551 -200
rect -5873 -4331 -5551 -4330
rect -6296 -4678 -6192 -4382
rect -6885 -4730 -6563 -4729
rect -6885 -8860 -6884 -4730
rect -6564 -8860 -6563 -4730
rect -6885 -8861 -6563 -8860
rect -7308 -9208 -7204 -8912
rect -7897 -9260 -7575 -9259
rect -7897 -13390 -7896 -9260
rect -7576 -13390 -7575 -9260
rect -7897 -13391 -7575 -13390
rect -7788 -13789 -7684 -13391
rect -7308 -13442 -7288 -9208
rect -7224 -13442 -7204 -9208
rect -6776 -9259 -6672 -8861
rect -6296 -8912 -6276 -4678
rect -6212 -8912 -6192 -4678
rect -5764 -4729 -5660 -4331
rect -5284 -4382 -5264 -148
rect -5200 -4382 -5180 -148
rect -4752 -199 -4648 199
rect -4272 148 -4252 4382
rect -4188 148 -4168 4382
rect -3740 4331 -3636 4729
rect -3260 4678 -3240 8912
rect -3176 4678 -3156 8912
rect -2728 8861 -2624 9259
rect -2248 9208 -2228 13442
rect -2164 9208 -2144 13442
rect -1716 13391 -1612 13789
rect -1236 13738 -1216 17972
rect -1152 13738 -1132 17972
rect -704 17921 -600 18120
rect -224 17972 -120 18120
rect -813 17920 -491 17921
rect -813 13790 -812 17920
rect -492 13790 -491 17920
rect -813 13789 -491 13790
rect -1236 13442 -1132 13738
rect -1825 13390 -1503 13391
rect -1825 9260 -1824 13390
rect -1504 9260 -1503 13390
rect -1825 9259 -1503 9260
rect -2248 8912 -2144 9208
rect -2837 8860 -2515 8861
rect -2837 4730 -2836 8860
rect -2516 4730 -2515 8860
rect -2837 4729 -2515 4730
rect -3260 4382 -3156 4678
rect -3849 4330 -3527 4331
rect -3849 200 -3848 4330
rect -3528 200 -3527 4330
rect -3849 199 -3527 200
rect -4272 -148 -4168 148
rect -4861 -200 -4539 -199
rect -4861 -4330 -4860 -200
rect -4540 -4330 -4539 -200
rect -4861 -4331 -4539 -4330
rect -5284 -4678 -5180 -4382
rect -5873 -4730 -5551 -4729
rect -5873 -8860 -5872 -4730
rect -5552 -8860 -5551 -4730
rect -5873 -8861 -5551 -8860
rect -6296 -9208 -6192 -8912
rect -6885 -9260 -6563 -9259
rect -6885 -13390 -6884 -9260
rect -6564 -13390 -6563 -9260
rect -6885 -13391 -6563 -13390
rect -7308 -13738 -7204 -13442
rect -7897 -13790 -7575 -13789
rect -7897 -17920 -7896 -13790
rect -7576 -17920 -7575 -13790
rect -7897 -17921 -7575 -17920
rect -7788 -18120 -7684 -17921
rect -7308 -17972 -7288 -13738
rect -7224 -17972 -7204 -13738
rect -6776 -13789 -6672 -13391
rect -6296 -13442 -6276 -9208
rect -6212 -13442 -6192 -9208
rect -5764 -9259 -5660 -8861
rect -5284 -8912 -5264 -4678
rect -5200 -8912 -5180 -4678
rect -4752 -4729 -4648 -4331
rect -4272 -4382 -4252 -148
rect -4188 -4382 -4168 -148
rect -3740 -199 -3636 199
rect -3260 148 -3240 4382
rect -3176 148 -3156 4382
rect -2728 4331 -2624 4729
rect -2248 4678 -2228 8912
rect -2164 4678 -2144 8912
rect -1716 8861 -1612 9259
rect -1236 9208 -1216 13442
rect -1152 9208 -1132 13442
rect -704 13391 -600 13789
rect -224 13738 -204 17972
rect -140 13738 -120 17972
rect 308 17921 412 18120
rect 788 17972 892 18120
rect 199 17920 521 17921
rect 199 13790 200 17920
rect 520 13790 521 17920
rect 199 13789 521 13790
rect -224 13442 -120 13738
rect -813 13390 -491 13391
rect -813 9260 -812 13390
rect -492 9260 -491 13390
rect -813 9259 -491 9260
rect -1236 8912 -1132 9208
rect -1825 8860 -1503 8861
rect -1825 4730 -1824 8860
rect -1504 4730 -1503 8860
rect -1825 4729 -1503 4730
rect -2248 4382 -2144 4678
rect -2837 4330 -2515 4331
rect -2837 200 -2836 4330
rect -2516 200 -2515 4330
rect -2837 199 -2515 200
rect -3260 -148 -3156 148
rect -3849 -200 -3527 -199
rect -3849 -4330 -3848 -200
rect -3528 -4330 -3527 -200
rect -3849 -4331 -3527 -4330
rect -4272 -4678 -4168 -4382
rect -4861 -4730 -4539 -4729
rect -4861 -8860 -4860 -4730
rect -4540 -8860 -4539 -4730
rect -4861 -8861 -4539 -8860
rect -5284 -9208 -5180 -8912
rect -5873 -9260 -5551 -9259
rect -5873 -13390 -5872 -9260
rect -5552 -13390 -5551 -9260
rect -5873 -13391 -5551 -13390
rect -6296 -13738 -6192 -13442
rect -6885 -13790 -6563 -13789
rect -6885 -17920 -6884 -13790
rect -6564 -17920 -6563 -13790
rect -6885 -17921 -6563 -17920
rect -7308 -18120 -7204 -17972
rect -6776 -18120 -6672 -17921
rect -6296 -17972 -6276 -13738
rect -6212 -17972 -6192 -13738
rect -5764 -13789 -5660 -13391
rect -5284 -13442 -5264 -9208
rect -5200 -13442 -5180 -9208
rect -4752 -9259 -4648 -8861
rect -4272 -8912 -4252 -4678
rect -4188 -8912 -4168 -4678
rect -3740 -4729 -3636 -4331
rect -3260 -4382 -3240 -148
rect -3176 -4382 -3156 -148
rect -2728 -199 -2624 199
rect -2248 148 -2228 4382
rect -2164 148 -2144 4382
rect -1716 4331 -1612 4729
rect -1236 4678 -1216 8912
rect -1152 4678 -1132 8912
rect -704 8861 -600 9259
rect -224 9208 -204 13442
rect -140 9208 -120 13442
rect 308 13391 412 13789
rect 788 13738 808 17972
rect 872 13738 892 17972
rect 1320 17921 1424 18120
rect 1800 17972 1904 18120
rect 1211 17920 1533 17921
rect 1211 13790 1212 17920
rect 1532 13790 1533 17920
rect 1211 13789 1533 13790
rect 788 13442 892 13738
rect 199 13390 521 13391
rect 199 9260 200 13390
rect 520 9260 521 13390
rect 199 9259 521 9260
rect -224 8912 -120 9208
rect -813 8860 -491 8861
rect -813 4730 -812 8860
rect -492 4730 -491 8860
rect -813 4729 -491 4730
rect -1236 4382 -1132 4678
rect -1825 4330 -1503 4331
rect -1825 200 -1824 4330
rect -1504 200 -1503 4330
rect -1825 199 -1503 200
rect -2248 -148 -2144 148
rect -2837 -200 -2515 -199
rect -2837 -4330 -2836 -200
rect -2516 -4330 -2515 -200
rect -2837 -4331 -2515 -4330
rect -3260 -4678 -3156 -4382
rect -3849 -4730 -3527 -4729
rect -3849 -8860 -3848 -4730
rect -3528 -8860 -3527 -4730
rect -3849 -8861 -3527 -8860
rect -4272 -9208 -4168 -8912
rect -4861 -9260 -4539 -9259
rect -4861 -13390 -4860 -9260
rect -4540 -13390 -4539 -9260
rect -4861 -13391 -4539 -13390
rect -5284 -13738 -5180 -13442
rect -5873 -13790 -5551 -13789
rect -5873 -17920 -5872 -13790
rect -5552 -17920 -5551 -13790
rect -5873 -17921 -5551 -17920
rect -6296 -18120 -6192 -17972
rect -5764 -18120 -5660 -17921
rect -5284 -17972 -5264 -13738
rect -5200 -17972 -5180 -13738
rect -4752 -13789 -4648 -13391
rect -4272 -13442 -4252 -9208
rect -4188 -13442 -4168 -9208
rect -3740 -9259 -3636 -8861
rect -3260 -8912 -3240 -4678
rect -3176 -8912 -3156 -4678
rect -2728 -4729 -2624 -4331
rect -2248 -4382 -2228 -148
rect -2164 -4382 -2144 -148
rect -1716 -199 -1612 199
rect -1236 148 -1216 4382
rect -1152 148 -1132 4382
rect -704 4331 -600 4729
rect -224 4678 -204 8912
rect -140 4678 -120 8912
rect 308 8861 412 9259
rect 788 9208 808 13442
rect 872 9208 892 13442
rect 1320 13391 1424 13789
rect 1800 13738 1820 17972
rect 1884 13738 1904 17972
rect 2332 17921 2436 18120
rect 2812 17972 2916 18120
rect 2223 17920 2545 17921
rect 2223 13790 2224 17920
rect 2544 13790 2545 17920
rect 2223 13789 2545 13790
rect 1800 13442 1904 13738
rect 1211 13390 1533 13391
rect 1211 9260 1212 13390
rect 1532 9260 1533 13390
rect 1211 9259 1533 9260
rect 788 8912 892 9208
rect 199 8860 521 8861
rect 199 4730 200 8860
rect 520 4730 521 8860
rect 199 4729 521 4730
rect -224 4382 -120 4678
rect -813 4330 -491 4331
rect -813 200 -812 4330
rect -492 200 -491 4330
rect -813 199 -491 200
rect -1236 -148 -1132 148
rect -1825 -200 -1503 -199
rect -1825 -4330 -1824 -200
rect -1504 -4330 -1503 -200
rect -1825 -4331 -1503 -4330
rect -2248 -4678 -2144 -4382
rect -2837 -4730 -2515 -4729
rect -2837 -8860 -2836 -4730
rect -2516 -8860 -2515 -4730
rect -2837 -8861 -2515 -8860
rect -3260 -9208 -3156 -8912
rect -3849 -9260 -3527 -9259
rect -3849 -13390 -3848 -9260
rect -3528 -13390 -3527 -9260
rect -3849 -13391 -3527 -13390
rect -4272 -13738 -4168 -13442
rect -4861 -13790 -4539 -13789
rect -4861 -17920 -4860 -13790
rect -4540 -17920 -4539 -13790
rect -4861 -17921 -4539 -17920
rect -5284 -18120 -5180 -17972
rect -4752 -18120 -4648 -17921
rect -4272 -17972 -4252 -13738
rect -4188 -17972 -4168 -13738
rect -3740 -13789 -3636 -13391
rect -3260 -13442 -3240 -9208
rect -3176 -13442 -3156 -9208
rect -2728 -9259 -2624 -8861
rect -2248 -8912 -2228 -4678
rect -2164 -8912 -2144 -4678
rect -1716 -4729 -1612 -4331
rect -1236 -4382 -1216 -148
rect -1152 -4382 -1132 -148
rect -704 -199 -600 199
rect -224 148 -204 4382
rect -140 148 -120 4382
rect 308 4331 412 4729
rect 788 4678 808 8912
rect 872 4678 892 8912
rect 1320 8861 1424 9259
rect 1800 9208 1820 13442
rect 1884 9208 1904 13442
rect 2332 13391 2436 13789
rect 2812 13738 2832 17972
rect 2896 13738 2916 17972
rect 3344 17921 3448 18120
rect 3824 17972 3928 18120
rect 3235 17920 3557 17921
rect 3235 13790 3236 17920
rect 3556 13790 3557 17920
rect 3235 13789 3557 13790
rect 2812 13442 2916 13738
rect 2223 13390 2545 13391
rect 2223 9260 2224 13390
rect 2544 9260 2545 13390
rect 2223 9259 2545 9260
rect 1800 8912 1904 9208
rect 1211 8860 1533 8861
rect 1211 4730 1212 8860
rect 1532 4730 1533 8860
rect 1211 4729 1533 4730
rect 788 4382 892 4678
rect 199 4330 521 4331
rect 199 200 200 4330
rect 520 200 521 4330
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -4330 -812 -200
rect -492 -4330 -491 -200
rect -813 -4331 -491 -4330
rect -1236 -4678 -1132 -4382
rect -1825 -4730 -1503 -4729
rect -1825 -8860 -1824 -4730
rect -1504 -8860 -1503 -4730
rect -1825 -8861 -1503 -8860
rect -2248 -9208 -2144 -8912
rect -2837 -9260 -2515 -9259
rect -2837 -13390 -2836 -9260
rect -2516 -13390 -2515 -9260
rect -2837 -13391 -2515 -13390
rect -3260 -13738 -3156 -13442
rect -3849 -13790 -3527 -13789
rect -3849 -17920 -3848 -13790
rect -3528 -17920 -3527 -13790
rect -3849 -17921 -3527 -17920
rect -4272 -18120 -4168 -17972
rect -3740 -18120 -3636 -17921
rect -3260 -17972 -3240 -13738
rect -3176 -17972 -3156 -13738
rect -2728 -13789 -2624 -13391
rect -2248 -13442 -2228 -9208
rect -2164 -13442 -2144 -9208
rect -1716 -9259 -1612 -8861
rect -1236 -8912 -1216 -4678
rect -1152 -8912 -1132 -4678
rect -704 -4729 -600 -4331
rect -224 -4382 -204 -148
rect -140 -4382 -120 -148
rect 308 -199 412 199
rect 788 148 808 4382
rect 872 148 892 4382
rect 1320 4331 1424 4729
rect 1800 4678 1820 8912
rect 1884 4678 1904 8912
rect 2332 8861 2436 9259
rect 2812 9208 2832 13442
rect 2896 9208 2916 13442
rect 3344 13391 3448 13789
rect 3824 13738 3844 17972
rect 3908 13738 3928 17972
rect 4356 17921 4460 18120
rect 4836 17972 4940 18120
rect 4247 17920 4569 17921
rect 4247 13790 4248 17920
rect 4568 13790 4569 17920
rect 4247 13789 4569 13790
rect 3824 13442 3928 13738
rect 3235 13390 3557 13391
rect 3235 9260 3236 13390
rect 3556 9260 3557 13390
rect 3235 9259 3557 9260
rect 2812 8912 2916 9208
rect 2223 8860 2545 8861
rect 2223 4730 2224 8860
rect 2544 4730 2545 8860
rect 2223 4729 2545 4730
rect 1800 4382 1904 4678
rect 1211 4330 1533 4331
rect 1211 200 1212 4330
rect 1532 200 1533 4330
rect 1211 199 1533 200
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -4330 200 -200
rect 520 -4330 521 -200
rect 199 -4331 521 -4330
rect -224 -4678 -120 -4382
rect -813 -4730 -491 -4729
rect -813 -8860 -812 -4730
rect -492 -8860 -491 -4730
rect -813 -8861 -491 -8860
rect -1236 -9208 -1132 -8912
rect -1825 -9260 -1503 -9259
rect -1825 -13390 -1824 -9260
rect -1504 -13390 -1503 -9260
rect -1825 -13391 -1503 -13390
rect -2248 -13738 -2144 -13442
rect -2837 -13790 -2515 -13789
rect -2837 -17920 -2836 -13790
rect -2516 -17920 -2515 -13790
rect -2837 -17921 -2515 -17920
rect -3260 -18120 -3156 -17972
rect -2728 -18120 -2624 -17921
rect -2248 -17972 -2228 -13738
rect -2164 -17972 -2144 -13738
rect -1716 -13789 -1612 -13391
rect -1236 -13442 -1216 -9208
rect -1152 -13442 -1132 -9208
rect -704 -9259 -600 -8861
rect -224 -8912 -204 -4678
rect -140 -8912 -120 -4678
rect 308 -4729 412 -4331
rect 788 -4382 808 -148
rect 872 -4382 892 -148
rect 1320 -199 1424 199
rect 1800 148 1820 4382
rect 1884 148 1904 4382
rect 2332 4331 2436 4729
rect 2812 4678 2832 8912
rect 2896 4678 2916 8912
rect 3344 8861 3448 9259
rect 3824 9208 3844 13442
rect 3908 9208 3928 13442
rect 4356 13391 4460 13789
rect 4836 13738 4856 17972
rect 4920 13738 4940 17972
rect 5368 17921 5472 18120
rect 5848 17972 5952 18120
rect 5259 17920 5581 17921
rect 5259 13790 5260 17920
rect 5580 13790 5581 17920
rect 5259 13789 5581 13790
rect 4836 13442 4940 13738
rect 4247 13390 4569 13391
rect 4247 9260 4248 13390
rect 4568 9260 4569 13390
rect 4247 9259 4569 9260
rect 3824 8912 3928 9208
rect 3235 8860 3557 8861
rect 3235 4730 3236 8860
rect 3556 4730 3557 8860
rect 3235 4729 3557 4730
rect 2812 4382 2916 4678
rect 2223 4330 2545 4331
rect 2223 200 2224 4330
rect 2544 200 2545 4330
rect 2223 199 2545 200
rect 1800 -148 1904 148
rect 1211 -200 1533 -199
rect 1211 -4330 1212 -200
rect 1532 -4330 1533 -200
rect 1211 -4331 1533 -4330
rect 788 -4678 892 -4382
rect 199 -4730 521 -4729
rect 199 -8860 200 -4730
rect 520 -8860 521 -4730
rect 199 -8861 521 -8860
rect -224 -9208 -120 -8912
rect -813 -9260 -491 -9259
rect -813 -13390 -812 -9260
rect -492 -13390 -491 -9260
rect -813 -13391 -491 -13390
rect -1236 -13738 -1132 -13442
rect -1825 -13790 -1503 -13789
rect -1825 -17920 -1824 -13790
rect -1504 -17920 -1503 -13790
rect -1825 -17921 -1503 -17920
rect -2248 -18120 -2144 -17972
rect -1716 -18120 -1612 -17921
rect -1236 -17972 -1216 -13738
rect -1152 -17972 -1132 -13738
rect -704 -13789 -600 -13391
rect -224 -13442 -204 -9208
rect -140 -13442 -120 -9208
rect 308 -9259 412 -8861
rect 788 -8912 808 -4678
rect 872 -8912 892 -4678
rect 1320 -4729 1424 -4331
rect 1800 -4382 1820 -148
rect 1884 -4382 1904 -148
rect 2332 -199 2436 199
rect 2812 148 2832 4382
rect 2896 148 2916 4382
rect 3344 4331 3448 4729
rect 3824 4678 3844 8912
rect 3908 4678 3928 8912
rect 4356 8861 4460 9259
rect 4836 9208 4856 13442
rect 4920 9208 4940 13442
rect 5368 13391 5472 13789
rect 5848 13738 5868 17972
rect 5932 13738 5952 17972
rect 6380 17921 6484 18120
rect 6860 17972 6964 18120
rect 6271 17920 6593 17921
rect 6271 13790 6272 17920
rect 6592 13790 6593 17920
rect 6271 13789 6593 13790
rect 5848 13442 5952 13738
rect 5259 13390 5581 13391
rect 5259 9260 5260 13390
rect 5580 9260 5581 13390
rect 5259 9259 5581 9260
rect 4836 8912 4940 9208
rect 4247 8860 4569 8861
rect 4247 4730 4248 8860
rect 4568 4730 4569 8860
rect 4247 4729 4569 4730
rect 3824 4382 3928 4678
rect 3235 4330 3557 4331
rect 3235 200 3236 4330
rect 3556 200 3557 4330
rect 3235 199 3557 200
rect 2812 -148 2916 148
rect 2223 -200 2545 -199
rect 2223 -4330 2224 -200
rect 2544 -4330 2545 -200
rect 2223 -4331 2545 -4330
rect 1800 -4678 1904 -4382
rect 1211 -4730 1533 -4729
rect 1211 -8860 1212 -4730
rect 1532 -8860 1533 -4730
rect 1211 -8861 1533 -8860
rect 788 -9208 892 -8912
rect 199 -9260 521 -9259
rect 199 -13390 200 -9260
rect 520 -13390 521 -9260
rect 199 -13391 521 -13390
rect -224 -13738 -120 -13442
rect -813 -13790 -491 -13789
rect -813 -17920 -812 -13790
rect -492 -17920 -491 -13790
rect -813 -17921 -491 -17920
rect -1236 -18120 -1132 -17972
rect -704 -18120 -600 -17921
rect -224 -17972 -204 -13738
rect -140 -17972 -120 -13738
rect 308 -13789 412 -13391
rect 788 -13442 808 -9208
rect 872 -13442 892 -9208
rect 1320 -9259 1424 -8861
rect 1800 -8912 1820 -4678
rect 1884 -8912 1904 -4678
rect 2332 -4729 2436 -4331
rect 2812 -4382 2832 -148
rect 2896 -4382 2916 -148
rect 3344 -199 3448 199
rect 3824 148 3844 4382
rect 3908 148 3928 4382
rect 4356 4331 4460 4729
rect 4836 4678 4856 8912
rect 4920 4678 4940 8912
rect 5368 8861 5472 9259
rect 5848 9208 5868 13442
rect 5932 9208 5952 13442
rect 6380 13391 6484 13789
rect 6860 13738 6880 17972
rect 6944 13738 6964 17972
rect 7392 17921 7496 18120
rect 7872 17972 7976 18120
rect 7283 17920 7605 17921
rect 7283 13790 7284 17920
rect 7604 13790 7605 17920
rect 7283 13789 7605 13790
rect 6860 13442 6964 13738
rect 6271 13390 6593 13391
rect 6271 9260 6272 13390
rect 6592 9260 6593 13390
rect 6271 9259 6593 9260
rect 5848 8912 5952 9208
rect 5259 8860 5581 8861
rect 5259 4730 5260 8860
rect 5580 4730 5581 8860
rect 5259 4729 5581 4730
rect 4836 4382 4940 4678
rect 4247 4330 4569 4331
rect 4247 200 4248 4330
rect 4568 200 4569 4330
rect 4247 199 4569 200
rect 3824 -148 3928 148
rect 3235 -200 3557 -199
rect 3235 -4330 3236 -200
rect 3556 -4330 3557 -200
rect 3235 -4331 3557 -4330
rect 2812 -4678 2916 -4382
rect 2223 -4730 2545 -4729
rect 2223 -8860 2224 -4730
rect 2544 -8860 2545 -4730
rect 2223 -8861 2545 -8860
rect 1800 -9208 1904 -8912
rect 1211 -9260 1533 -9259
rect 1211 -13390 1212 -9260
rect 1532 -13390 1533 -9260
rect 1211 -13391 1533 -13390
rect 788 -13738 892 -13442
rect 199 -13790 521 -13789
rect 199 -17920 200 -13790
rect 520 -17920 521 -13790
rect 199 -17921 521 -17920
rect -224 -18120 -120 -17972
rect 308 -18120 412 -17921
rect 788 -17972 808 -13738
rect 872 -17972 892 -13738
rect 1320 -13789 1424 -13391
rect 1800 -13442 1820 -9208
rect 1884 -13442 1904 -9208
rect 2332 -9259 2436 -8861
rect 2812 -8912 2832 -4678
rect 2896 -8912 2916 -4678
rect 3344 -4729 3448 -4331
rect 3824 -4382 3844 -148
rect 3908 -4382 3928 -148
rect 4356 -199 4460 199
rect 4836 148 4856 4382
rect 4920 148 4940 4382
rect 5368 4331 5472 4729
rect 5848 4678 5868 8912
rect 5932 4678 5952 8912
rect 6380 8861 6484 9259
rect 6860 9208 6880 13442
rect 6944 9208 6964 13442
rect 7392 13391 7496 13789
rect 7872 13738 7892 17972
rect 7956 13738 7976 17972
rect 7872 13442 7976 13738
rect 7283 13390 7605 13391
rect 7283 9260 7284 13390
rect 7604 9260 7605 13390
rect 7283 9259 7605 9260
rect 6860 8912 6964 9208
rect 6271 8860 6593 8861
rect 6271 4730 6272 8860
rect 6592 4730 6593 8860
rect 6271 4729 6593 4730
rect 5848 4382 5952 4678
rect 5259 4330 5581 4331
rect 5259 200 5260 4330
rect 5580 200 5581 4330
rect 5259 199 5581 200
rect 4836 -148 4940 148
rect 4247 -200 4569 -199
rect 4247 -4330 4248 -200
rect 4568 -4330 4569 -200
rect 4247 -4331 4569 -4330
rect 3824 -4678 3928 -4382
rect 3235 -4730 3557 -4729
rect 3235 -8860 3236 -4730
rect 3556 -8860 3557 -4730
rect 3235 -8861 3557 -8860
rect 2812 -9208 2916 -8912
rect 2223 -9260 2545 -9259
rect 2223 -13390 2224 -9260
rect 2544 -13390 2545 -9260
rect 2223 -13391 2545 -13390
rect 1800 -13738 1904 -13442
rect 1211 -13790 1533 -13789
rect 1211 -17920 1212 -13790
rect 1532 -17920 1533 -13790
rect 1211 -17921 1533 -17920
rect 788 -18120 892 -17972
rect 1320 -18120 1424 -17921
rect 1800 -17972 1820 -13738
rect 1884 -17972 1904 -13738
rect 2332 -13789 2436 -13391
rect 2812 -13442 2832 -9208
rect 2896 -13442 2916 -9208
rect 3344 -9259 3448 -8861
rect 3824 -8912 3844 -4678
rect 3908 -8912 3928 -4678
rect 4356 -4729 4460 -4331
rect 4836 -4382 4856 -148
rect 4920 -4382 4940 -148
rect 5368 -199 5472 199
rect 5848 148 5868 4382
rect 5932 148 5952 4382
rect 6380 4331 6484 4729
rect 6860 4678 6880 8912
rect 6944 4678 6964 8912
rect 7392 8861 7496 9259
rect 7872 9208 7892 13442
rect 7956 9208 7976 13442
rect 7872 8912 7976 9208
rect 7283 8860 7605 8861
rect 7283 4730 7284 8860
rect 7604 4730 7605 8860
rect 7283 4729 7605 4730
rect 6860 4382 6964 4678
rect 6271 4330 6593 4331
rect 6271 200 6272 4330
rect 6592 200 6593 4330
rect 6271 199 6593 200
rect 5848 -148 5952 148
rect 5259 -200 5581 -199
rect 5259 -4330 5260 -200
rect 5580 -4330 5581 -200
rect 5259 -4331 5581 -4330
rect 4836 -4678 4940 -4382
rect 4247 -4730 4569 -4729
rect 4247 -8860 4248 -4730
rect 4568 -8860 4569 -4730
rect 4247 -8861 4569 -8860
rect 3824 -9208 3928 -8912
rect 3235 -9260 3557 -9259
rect 3235 -13390 3236 -9260
rect 3556 -13390 3557 -9260
rect 3235 -13391 3557 -13390
rect 2812 -13738 2916 -13442
rect 2223 -13790 2545 -13789
rect 2223 -17920 2224 -13790
rect 2544 -17920 2545 -13790
rect 2223 -17921 2545 -17920
rect 1800 -18120 1904 -17972
rect 2332 -18120 2436 -17921
rect 2812 -17972 2832 -13738
rect 2896 -17972 2916 -13738
rect 3344 -13789 3448 -13391
rect 3824 -13442 3844 -9208
rect 3908 -13442 3928 -9208
rect 4356 -9259 4460 -8861
rect 4836 -8912 4856 -4678
rect 4920 -8912 4940 -4678
rect 5368 -4729 5472 -4331
rect 5848 -4382 5868 -148
rect 5932 -4382 5952 -148
rect 6380 -199 6484 199
rect 6860 148 6880 4382
rect 6944 148 6964 4382
rect 7392 4331 7496 4729
rect 7872 4678 7892 8912
rect 7956 4678 7976 8912
rect 7872 4382 7976 4678
rect 7283 4330 7605 4331
rect 7283 200 7284 4330
rect 7604 200 7605 4330
rect 7283 199 7605 200
rect 6860 -148 6964 148
rect 6271 -200 6593 -199
rect 6271 -4330 6272 -200
rect 6592 -4330 6593 -200
rect 6271 -4331 6593 -4330
rect 5848 -4678 5952 -4382
rect 5259 -4730 5581 -4729
rect 5259 -8860 5260 -4730
rect 5580 -8860 5581 -4730
rect 5259 -8861 5581 -8860
rect 4836 -9208 4940 -8912
rect 4247 -9260 4569 -9259
rect 4247 -13390 4248 -9260
rect 4568 -13390 4569 -9260
rect 4247 -13391 4569 -13390
rect 3824 -13738 3928 -13442
rect 3235 -13790 3557 -13789
rect 3235 -17920 3236 -13790
rect 3556 -17920 3557 -13790
rect 3235 -17921 3557 -17920
rect 2812 -18120 2916 -17972
rect 3344 -18120 3448 -17921
rect 3824 -17972 3844 -13738
rect 3908 -17972 3928 -13738
rect 4356 -13789 4460 -13391
rect 4836 -13442 4856 -9208
rect 4920 -13442 4940 -9208
rect 5368 -9259 5472 -8861
rect 5848 -8912 5868 -4678
rect 5932 -8912 5952 -4678
rect 6380 -4729 6484 -4331
rect 6860 -4382 6880 -148
rect 6944 -4382 6964 -148
rect 7392 -199 7496 199
rect 7872 148 7892 4382
rect 7956 148 7976 4382
rect 7872 -148 7976 148
rect 7283 -200 7605 -199
rect 7283 -4330 7284 -200
rect 7604 -4330 7605 -200
rect 7283 -4331 7605 -4330
rect 6860 -4678 6964 -4382
rect 6271 -4730 6593 -4729
rect 6271 -8860 6272 -4730
rect 6592 -8860 6593 -4730
rect 6271 -8861 6593 -8860
rect 5848 -9208 5952 -8912
rect 5259 -9260 5581 -9259
rect 5259 -13390 5260 -9260
rect 5580 -13390 5581 -9260
rect 5259 -13391 5581 -13390
rect 4836 -13738 4940 -13442
rect 4247 -13790 4569 -13789
rect 4247 -17920 4248 -13790
rect 4568 -17920 4569 -13790
rect 4247 -17921 4569 -17920
rect 3824 -18120 3928 -17972
rect 4356 -18120 4460 -17921
rect 4836 -17972 4856 -13738
rect 4920 -17972 4940 -13738
rect 5368 -13789 5472 -13391
rect 5848 -13442 5868 -9208
rect 5932 -13442 5952 -9208
rect 6380 -9259 6484 -8861
rect 6860 -8912 6880 -4678
rect 6944 -8912 6964 -4678
rect 7392 -4729 7496 -4331
rect 7872 -4382 7892 -148
rect 7956 -4382 7976 -148
rect 7872 -4678 7976 -4382
rect 7283 -4730 7605 -4729
rect 7283 -8860 7284 -4730
rect 7604 -8860 7605 -4730
rect 7283 -8861 7605 -8860
rect 6860 -9208 6964 -8912
rect 6271 -9260 6593 -9259
rect 6271 -13390 6272 -9260
rect 6592 -13390 6593 -9260
rect 6271 -13391 6593 -13390
rect 5848 -13738 5952 -13442
rect 5259 -13790 5581 -13789
rect 5259 -17920 5260 -13790
rect 5580 -17920 5581 -13790
rect 5259 -17921 5581 -17920
rect 4836 -18120 4940 -17972
rect 5368 -18120 5472 -17921
rect 5848 -17972 5868 -13738
rect 5932 -17972 5952 -13738
rect 6380 -13789 6484 -13391
rect 6860 -13442 6880 -9208
rect 6944 -13442 6964 -9208
rect 7392 -9259 7496 -8861
rect 7872 -8912 7892 -4678
rect 7956 -8912 7976 -4678
rect 7872 -9208 7976 -8912
rect 7283 -9260 7605 -9259
rect 7283 -13390 7284 -9260
rect 7604 -13390 7605 -9260
rect 7283 -13391 7605 -13390
rect 6860 -13738 6964 -13442
rect 6271 -13790 6593 -13789
rect 6271 -17920 6272 -13790
rect 6592 -17920 6593 -13790
rect 6271 -17921 6593 -17920
rect 5848 -18120 5952 -17972
rect 6380 -18120 6484 -17921
rect 6860 -17972 6880 -13738
rect 6944 -17972 6964 -13738
rect 7392 -13789 7496 -13391
rect 7872 -13442 7892 -9208
rect 7956 -13442 7976 -9208
rect 7872 -13738 7976 -13442
rect 7283 -13790 7605 -13789
rect 7283 -17920 7284 -13790
rect 7604 -17920 7605 -13790
rect 7283 -17921 7605 -17920
rect 6860 -18120 6964 -17972
rect 7392 -18120 7496 -17921
rect 7872 -17972 7892 -13738
rect 7956 -17972 7976 -13738
rect 7872 -18120 7976 -17972
<< properties >>
string FIXED_BBOX 7204 13710 7684 18000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 16 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
