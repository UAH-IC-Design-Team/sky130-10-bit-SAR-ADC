magic
tech sky130A
magscale 1 2
timestamp 1668286574
<< viali >>
rect 2053 21641 2087 21675
rect 3249 21641 3283 21675
rect 4629 21641 4663 21675
rect 5917 21641 5951 21675
rect 7297 21641 7331 21675
rect 8493 21641 8527 21675
rect 9873 21641 9907 21675
rect 10977 21641 11011 21675
rect 12357 21641 12391 21675
rect 14473 21641 14507 21675
rect 15209 21641 15243 21675
rect 17049 21641 17083 21675
rect 17785 21641 17819 21675
rect 19625 21641 19659 21675
rect 2237 21505 2271 21539
rect 3433 21505 3467 21539
rect 4813 21505 4847 21539
rect 5733 21505 5767 21539
rect 7113 21505 7147 21539
rect 8309 21505 8343 21539
rect 9689 21505 9723 21539
rect 11161 21505 11195 21539
rect 12541 21505 12575 21539
rect 14289 21505 14323 21539
rect 15025 21505 15059 21539
rect 15910 21505 15944 21539
rect 16865 21505 16899 21539
rect 17601 21505 17635 21539
rect 18889 21505 18923 21539
rect 19441 21505 19475 21539
rect 18705 21369 18739 21403
rect 15807 21301 15841 21335
rect 1777 21097 1811 21131
rect 17187 21097 17221 21131
rect 20085 21097 20119 21131
rect 6285 20961 6319 20995
rect 13737 20961 13771 20995
rect 15761 20961 15795 20995
rect 1593 20893 1627 20927
rect 2697 20893 2731 20927
rect 6561 20893 6595 20927
rect 7021 20893 7055 20927
rect 7205 20893 7239 20927
rect 8192 20893 8226 20927
rect 10149 20893 10183 20927
rect 13461 20893 13495 20927
rect 15393 20893 15427 20927
rect 17842 20893 17876 20927
rect 18454 20893 18488 20927
rect 19901 20893 19935 20927
rect 3249 20825 3283 20859
rect 10425 20825 10459 20859
rect 4813 20757 4847 20791
rect 8263 20757 8297 20791
rect 11897 20757 11931 20791
rect 17739 20757 17773 20791
rect 18383 20757 18417 20791
rect 1685 20553 1719 20587
rect 9735 20553 9769 20587
rect 13553 20553 13587 20587
rect 18659 20553 18693 20587
rect 19257 20553 19291 20587
rect 4721 20485 4755 20519
rect 5871 20485 5905 20519
rect 14289 20485 14323 20519
rect 1869 20417 1903 20451
rect 2605 20417 2639 20451
rect 5974 20417 6008 20451
rect 7389 20417 7423 20451
rect 8309 20417 8343 20451
rect 11805 20417 11839 20451
rect 17233 20417 17267 20451
rect 19441 20417 19475 20451
rect 19901 20417 19935 20451
rect 3249 20349 3283 20383
rect 4997 20349 5031 20383
rect 7941 20349 7975 20383
rect 12081 20349 12115 20383
rect 14013 20349 14047 20383
rect 16865 20349 16899 20383
rect 2789 20213 2823 20247
rect 7113 20213 7147 20247
rect 15761 20213 15795 20247
rect 20085 20213 20119 20247
rect 2605 20009 2639 20043
rect 7757 20009 7791 20043
rect 12817 20009 12851 20043
rect 14289 20009 14323 20043
rect 18889 20009 18923 20043
rect 6285 19873 6319 19907
rect 11069 19873 11103 19907
rect 11345 19873 11379 19907
rect 15761 19873 15795 19907
rect 16037 19873 16071 19907
rect 17417 19873 17451 19907
rect 19441 19873 19475 19907
rect 2789 19805 2823 19839
rect 6009 19805 6043 19839
rect 16497 19805 16531 19839
rect 17141 19805 17175 19839
rect 19625 19805 19659 19839
rect 19809 19737 19843 19771
rect 16681 19669 16715 19703
rect 7021 19465 7055 19499
rect 10977 19465 11011 19499
rect 17647 19465 17681 19499
rect 2605 19397 2639 19431
rect 9505 19397 9539 19431
rect 8769 19329 8803 19363
rect 9229 19329 9263 19363
rect 16900 19329 16934 19363
rect 17576 19329 17610 19363
rect 2329 19261 2363 19295
rect 8493 19261 8527 19295
rect 18245 19261 18279 19295
rect 18521 19261 18555 19295
rect 4077 19125 4111 19159
rect 17003 19125 17037 19159
rect 19993 19125 20027 19159
rect 8585 18921 8619 18955
rect 12495 18921 12529 18955
rect 17877 18921 17911 18955
rect 3985 18785 4019 18819
rect 4261 18785 4295 18819
rect 11069 18785 11103 18819
rect 17509 18785 17543 18819
rect 6837 18717 6871 18751
rect 10701 18717 10735 18751
rect 15301 18717 15335 18751
rect 15945 18717 15979 18751
rect 16405 18717 16439 18751
rect 17049 18717 17083 18751
rect 17693 18717 17727 18751
rect 18486 18717 18520 18751
rect 20177 18717 20211 18751
rect 7113 18649 7147 18683
rect 5733 18581 5767 18615
rect 18383 18581 18417 18615
rect 19993 18581 20027 18615
rect 8309 18377 8343 18411
rect 11115 18377 11149 18411
rect 12495 18377 12529 18411
rect 16221 18377 16255 18411
rect 19625 18377 19659 18411
rect 5641 18309 5675 18343
rect 18153 18309 18187 18343
rect 2513 18241 2547 18275
rect 9321 18241 9355 18275
rect 11989 18241 12023 18275
rect 12566 18241 12600 18275
rect 14473 18241 14507 18275
rect 17049 18241 17083 18275
rect 5917 18173 5951 18207
rect 6561 18173 6595 18207
rect 6837 18173 6871 18207
rect 9689 18173 9723 18207
rect 14749 18173 14783 18207
rect 17233 18173 17267 18207
rect 17877 18173 17911 18207
rect 1869 18037 1903 18071
rect 4169 18037 4203 18071
rect 11805 18037 11839 18071
rect 16865 18037 16899 18071
rect 6837 17833 6871 17867
rect 9643 17833 9677 17867
rect 14841 17833 14875 17867
rect 17095 17833 17129 17867
rect 5365 17697 5399 17731
rect 11989 17697 12023 17731
rect 14381 17697 14415 17731
rect 17601 17697 17635 17731
rect 17785 17697 17819 17731
rect 1961 17629 1995 17663
rect 3214 17629 3248 17663
rect 5089 17629 5123 17663
rect 9540 17629 9574 17663
rect 11713 17629 11747 17663
rect 13737 17629 13771 17663
rect 14473 17629 14507 17663
rect 17024 17629 17058 17663
rect 18705 17629 18739 17663
rect 18889 17629 18923 17663
rect 10517 17561 10551 17595
rect 10701 17561 10735 17595
rect 19901 17561 19935 17595
rect 20085 17561 20119 17595
rect 2605 17493 2639 17527
rect 3111 17493 3145 17527
rect 7573 17493 7607 17527
rect 17969 17493 18003 17527
rect 1593 17289 1627 17323
rect 9689 17289 9723 17323
rect 12725 17289 12759 17323
rect 17003 17289 17037 17323
rect 3065 17221 3099 17255
rect 3341 17153 3375 17187
rect 3868 17153 3902 17187
rect 7297 17153 7331 17187
rect 7941 17153 7975 17187
rect 9505 17153 9539 17187
rect 12541 17153 12575 17187
rect 14657 17153 14691 17187
rect 16129 17153 16163 17187
rect 16900 17153 16934 17187
rect 17877 17153 17911 17187
rect 15301 17085 15335 17119
rect 15945 17085 15979 17119
rect 18153 17085 18187 17119
rect 15761 17017 15795 17051
rect 3939 16949 3973 16983
rect 7113 16949 7147 16983
rect 7757 16949 7791 16983
rect 19625 16949 19659 16983
rect 8585 16745 8619 16779
rect 12449 16745 12483 16779
rect 16037 16745 16071 16779
rect 3019 16677 3053 16711
rect 2145 16609 2179 16643
rect 2513 16609 2547 16643
rect 3985 16609 4019 16643
rect 6837 16609 6871 16643
rect 7113 16609 7147 16643
rect 10333 16609 10367 16643
rect 13461 16609 13495 16643
rect 13737 16609 13771 16643
rect 14565 16609 14599 16643
rect 16497 16609 16531 16643
rect 16773 16609 16807 16643
rect 2329 16541 2363 16575
rect 3122 16541 3156 16575
rect 4169 16541 4203 16575
rect 4353 16541 4387 16575
rect 4813 16541 4847 16575
rect 10057 16541 10091 16575
rect 12265 16541 12299 16575
rect 13369 16541 13403 16575
rect 14289 16541 14323 16575
rect 20177 16541 20211 16575
rect 4997 16405 5031 16439
rect 11805 16405 11839 16439
rect 18245 16405 18279 16439
rect 19993 16405 20027 16439
rect 3387 16201 3421 16235
rect 7205 16201 7239 16235
rect 10609 16201 10643 16235
rect 14565 16201 14599 16235
rect 15301 16201 15335 16235
rect 20177 16201 20211 16235
rect 8677 16133 8711 16167
rect 17141 16133 17175 16167
rect 1593 16065 1627 16099
rect 7021 16065 7055 16099
rect 7665 16065 7699 16099
rect 10793 16065 10827 16099
rect 12173 16065 12207 16099
rect 12817 16065 12851 16099
rect 13921 16065 13955 16099
rect 15485 16065 15519 16099
rect 16246 16065 16280 16099
rect 16957 16065 16991 16099
rect 1961 15997 1995 16031
rect 8401 15997 8435 16031
rect 10149 15997 10183 16031
rect 18429 15997 18463 16031
rect 18705 15997 18739 16031
rect 7849 15929 7883 15963
rect 12357 15929 12391 15963
rect 13001 15929 13035 15963
rect 15669 15929 15703 15963
rect 16175 15929 16209 15963
rect 1915 15657 1949 15691
rect 17325 15657 17359 15691
rect 7665 15589 7699 15623
rect 10057 15589 10091 15623
rect 18337 15589 18371 15623
rect 10609 15521 10643 15555
rect 10885 15521 10919 15555
rect 15117 15521 15151 15555
rect 2018 15453 2052 15487
rect 7481 15453 7515 15487
rect 9873 15453 9907 15487
rect 20085 15453 20119 15487
rect 15393 15385 15427 15419
rect 19717 15385 19751 15419
rect 12357 15317 12391 15351
rect 16865 15317 16899 15351
rect 18705 15317 18739 15351
rect 20177 15113 20211 15147
rect 18705 15045 18739 15079
rect 1593 14977 1627 15011
rect 5365 14977 5399 15011
rect 6929 14977 6963 15011
rect 7481 14977 7515 15011
rect 9229 14977 9263 15011
rect 10400 14977 10434 15011
rect 11989 14977 12023 15011
rect 14080 14977 14114 15011
rect 18429 14909 18463 14943
rect 7665 14841 7699 14875
rect 1777 14773 1811 14807
rect 5549 14773 5583 14807
rect 6837 14773 6871 14807
rect 9873 14773 9907 14807
rect 10471 14773 10505 14807
rect 12173 14773 12207 14807
rect 14151 14773 14185 14807
rect 10885 14569 10919 14603
rect 13093 14569 13127 14603
rect 16037 14569 16071 14603
rect 17049 14569 17083 14603
rect 4905 14501 4939 14535
rect 7941 14501 7975 14535
rect 11345 14501 11379 14535
rect 18061 14501 18095 14535
rect 5365 14433 5399 14467
rect 5641 14433 5675 14467
rect 9137 14433 9171 14467
rect 11529 14433 11563 14467
rect 14565 14433 14599 14467
rect 1685 14365 1719 14399
rect 4721 14365 4755 14399
rect 7757 14365 7791 14399
rect 12265 14365 12299 14399
rect 12909 14365 12943 14399
rect 14289 14365 14323 14399
rect 2789 14297 2823 14331
rect 9413 14297 9447 14331
rect 12449 14297 12483 14331
rect 1869 14229 1903 14263
rect 2697 14229 2731 14263
rect 7113 14229 7147 14263
rect 11713 14229 11747 14263
rect 18429 14229 18463 14263
rect 4031 14025 4065 14059
rect 4537 14025 4571 14059
rect 5549 14025 5583 14059
rect 7389 14025 7423 14059
rect 10609 14025 10643 14059
rect 14289 14025 14323 14059
rect 18705 13957 18739 13991
rect 1628 13889 1662 13923
rect 1731 13889 1765 13923
rect 2605 13889 2639 13923
rect 4721 13889 4755 13923
rect 5733 13889 5767 13923
rect 7205 13889 7239 13923
rect 8401 13889 8435 13923
rect 9965 13889 9999 13923
rect 11748 13889 11782 13923
rect 12541 13889 12575 13923
rect 2237 13821 2271 13855
rect 8309 13821 8343 13855
rect 8769 13821 8803 13855
rect 11851 13821 11885 13855
rect 12817 13821 12851 13855
rect 18429 13821 18463 13855
rect 20177 13685 20211 13719
rect 2145 13481 2179 13515
rect 11069 13481 11103 13515
rect 13323 13481 13357 13515
rect 14546 13481 14580 13515
rect 19993 13481 20027 13515
rect 2697 13413 2731 13447
rect 10701 13413 10735 13447
rect 12449 13413 12483 13447
rect 5549 13345 5583 13379
rect 5825 13345 5859 13379
rect 10885 13345 10919 13379
rect 12817 13345 12851 13379
rect 16773 13345 16807 13379
rect 1961 13277 1995 13311
rect 2881 13277 2915 13311
rect 12633 13277 12667 13311
rect 13426 13277 13460 13311
rect 14289 13277 14323 13311
rect 16497 13277 16531 13311
rect 20177 13277 20211 13311
rect 7297 13141 7331 13175
rect 16037 13141 16071 13175
rect 18245 13141 18279 13175
rect 2145 12937 2179 12971
rect 12725 12937 12759 12971
rect 16129 12937 16163 12971
rect 6837 12869 6871 12903
rect 15025 12869 15059 12903
rect 1961 12801 1995 12835
rect 2789 12801 2823 12835
rect 4353 12801 4387 12835
rect 8769 12801 8803 12835
rect 9965 12801 9999 12835
rect 12081 12801 12115 12835
rect 13670 12801 13704 12835
rect 16221 12801 16255 12835
rect 17417 12801 17451 12835
rect 6561 12733 6595 12767
rect 11897 12733 11931 12767
rect 12909 12733 12943 12767
rect 15301 12733 15335 12767
rect 17693 12733 17727 12767
rect 18429 12733 18463 12767
rect 18705 12733 18739 12767
rect 11713 12665 11747 12699
rect 13093 12665 13127 12699
rect 13599 12665 13633 12699
rect 2605 12597 2639 12631
rect 4537 12597 4571 12631
rect 8309 12597 8343 12631
rect 8953 12597 8987 12631
rect 10609 12597 10643 12631
rect 20177 12597 20211 12631
rect 6009 12393 6043 12427
rect 7573 12393 7607 12427
rect 10885 12393 10919 12427
rect 13461 12393 13495 12427
rect 17417 12393 17451 12427
rect 18797 12393 18831 12427
rect 8585 12325 8619 12359
rect 18429 12325 18463 12359
rect 19993 12325 20027 12359
rect 8125 12257 8159 12291
rect 9137 12257 9171 12291
rect 9413 12257 9447 12291
rect 15209 12257 15243 12291
rect 15485 12257 15519 12291
rect 1593 12189 1627 12223
rect 4721 12189 4755 12223
rect 5181 12189 5215 12223
rect 5825 12189 5859 12223
rect 6653 12189 6687 12223
rect 7389 12189 7423 12223
rect 8217 12189 8251 12223
rect 11713 12189 11747 12223
rect 14565 12189 14599 12223
rect 20177 12189 20211 12223
rect 11989 12121 12023 12155
rect 1777 12053 1811 12087
rect 4537 12053 4571 12087
rect 5365 12053 5399 12087
rect 6469 12053 6503 12087
rect 14381 12053 14415 12087
rect 16957 12053 16991 12087
rect 3709 11849 3743 11883
rect 4813 11849 4847 11883
rect 6653 11849 6687 11883
rect 11161 11849 11195 11883
rect 11943 11849 11977 11883
rect 16957 11849 16991 11883
rect 3525 11713 3559 11747
rect 4169 11713 4203 11747
rect 5825 11713 5859 11747
rect 6745 11713 6779 11747
rect 9940 11713 9974 11747
rect 10517 11713 10551 11747
rect 11872 11713 11906 11747
rect 13645 11713 13679 11747
rect 13921 11645 13955 11679
rect 15669 11645 15703 11679
rect 17969 11577 18003 11611
rect 6009 11509 6043 11543
rect 10011 11509 10045 11543
rect 18337 11509 18371 11543
rect 4629 11305 4663 11339
rect 5457 11305 5491 11339
rect 15209 11305 15243 11339
rect 15853 11305 15887 11339
rect 17693 11305 17727 11339
rect 1593 11237 1627 11271
rect 10425 11237 10459 11271
rect 16865 11237 16899 11271
rect 6193 11169 6227 11203
rect 6469 11169 6503 11203
rect 7941 11169 7975 11203
rect 10609 11169 10643 11203
rect 1777 11101 1811 11135
rect 3985 11101 4019 11135
rect 5273 11101 5307 11135
rect 8585 11101 8619 11135
rect 11412 11101 11446 11135
rect 17877 11101 17911 11135
rect 10793 11033 10827 11067
rect 14933 11033 14967 11067
rect 8401 10965 8435 10999
rect 11483 10965 11517 10999
rect 17233 10965 17267 10999
rect 3985 10761 4019 10795
rect 17969 10761 18003 10795
rect 10793 10693 10827 10727
rect 18705 10693 18739 10727
rect 1593 10625 1627 10659
rect 2237 10625 2271 10659
rect 3341 10625 3375 10659
rect 7757 10625 7791 10659
rect 8585 10625 8619 10659
rect 10977 10625 11011 10659
rect 13921 10625 13955 10659
rect 17785 10625 17819 10659
rect 7665 10557 7699 10591
rect 8861 10557 8895 10591
rect 11713 10557 11747 10591
rect 11989 10557 12023 10591
rect 14197 10557 14231 10591
rect 18429 10557 18463 10591
rect 8125 10489 8159 10523
rect 1777 10421 1811 10455
rect 2881 10421 2915 10455
rect 10333 10421 10367 10455
rect 13461 10421 13495 10455
rect 15669 10421 15703 10455
rect 20177 10421 20211 10455
rect 2329 10217 2363 10251
rect 3433 10217 3467 10251
rect 11437 10217 11471 10251
rect 12265 10217 12299 10251
rect 16037 10217 16071 10251
rect 19993 10217 20027 10251
rect 11897 10149 11931 10183
rect 11069 10081 11103 10115
rect 12081 10081 12115 10115
rect 1685 10013 1719 10047
rect 2789 10013 2823 10047
rect 8125 10013 8159 10047
rect 9388 10013 9422 10047
rect 9965 10013 9999 10047
rect 10609 10013 10643 10047
rect 11253 10013 11287 10047
rect 14289 10013 14323 10047
rect 20177 10013 20211 10047
rect 14565 9945 14599 9979
rect 8309 9877 8343 9911
rect 9459 9877 9493 9911
rect 9965 9673 9999 9707
rect 17785 9673 17819 9707
rect 4767 9605 4801 9639
rect 6837 9605 6871 9639
rect 18705 9605 18739 9639
rect 2053 9537 2087 9571
rect 9321 9537 9355 9571
rect 10609 9537 10643 9571
rect 10701 9537 10735 9571
rect 17969 9537 18003 9571
rect 1685 9469 1719 9503
rect 1961 9469 1995 9503
rect 2973 9469 3007 9503
rect 3341 9469 3375 9503
rect 18429 9469 18463 9503
rect 6929 9333 6963 9367
rect 10425 9333 10459 9367
rect 20177 9333 20211 9367
rect 3295 9129 3329 9163
rect 6837 9129 6871 9163
rect 18061 9129 18095 9163
rect 12725 9061 12759 9095
rect 19441 9061 19475 9095
rect 15393 8993 15427 9027
rect 16865 8993 16899 9027
rect 3398 8925 3432 8959
rect 4537 8925 4571 8959
rect 5089 8925 5123 8959
rect 7297 8925 7331 8959
rect 8125 8925 8159 8959
rect 9873 8925 9907 8959
rect 12541 8925 12575 8959
rect 13461 8925 13495 8959
rect 15117 8925 15151 8959
rect 17325 8925 17359 8959
rect 18245 8925 18279 8959
rect 18429 8925 18463 8959
rect 5365 8857 5399 8891
rect 19625 8857 19659 8891
rect 4353 8789 4387 8823
rect 7481 8789 7515 8823
rect 7941 8789 7975 8823
rect 9689 8789 9723 8823
rect 13277 8789 13311 8823
rect 17509 8789 17543 8823
rect 2513 8585 2547 8619
rect 5733 8585 5767 8619
rect 12081 8585 12115 8619
rect 15393 8585 15427 8619
rect 19993 8585 20027 8619
rect 6745 8517 6779 8551
rect 8401 8517 8435 8551
rect 17141 8517 17175 8551
rect 3985 8449 4019 8483
rect 7481 8449 7515 8483
rect 10333 8449 10367 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 14749 8449 14783 8483
rect 15577 8449 15611 8483
rect 16037 8449 16071 8483
rect 19257 8449 19291 8483
rect 20177 8449 20211 8483
rect 2697 8381 2731 8415
rect 4261 8381 4295 8415
rect 8125 8381 8159 8415
rect 12817 8381 12851 8415
rect 16865 8381 16899 8415
rect 2881 8313 2915 8347
rect 6561 8313 6595 8347
rect 7665 8313 7699 8347
rect 14933 8313 14967 8347
rect 16221 8313 16255 8347
rect 9873 8245 9907 8279
rect 10517 8245 10551 8279
rect 14289 8245 14323 8279
rect 18613 8245 18647 8279
rect 19073 8245 19107 8279
rect 4215 8041 4249 8075
rect 8585 8041 8619 8075
rect 9873 8041 9907 8075
rect 10964 8041 10998 8075
rect 12449 8041 12483 8075
rect 13093 8041 13127 8075
rect 16037 8041 16071 8075
rect 17325 8041 17359 8075
rect 3065 7973 3099 8007
rect 13737 7973 13771 8007
rect 16681 7973 16715 8007
rect 18429 7973 18463 8007
rect 19441 7973 19475 8007
rect 5319 7905 5353 7939
rect 7113 7905 7147 7939
rect 10701 7905 10735 7939
rect 14289 7905 14323 7939
rect 14565 7905 14599 7939
rect 18153 7905 18187 7939
rect 1777 7837 1811 7871
rect 3249 7837 3283 7871
rect 4318 7837 4352 7871
rect 5232 7837 5266 7871
rect 6837 7837 6871 7871
rect 9689 7837 9723 7871
rect 12909 7837 12943 7871
rect 13553 7837 13587 7871
rect 16497 7837 16531 7871
rect 17141 7837 17175 7871
rect 18061 7837 18095 7871
rect 19625 7837 19659 7871
rect 2421 7701 2455 7735
rect 3433 7701 3467 7735
rect 7205 7497 7239 7531
rect 11161 7497 11195 7531
rect 17969 7497 18003 7531
rect 9689 7429 9723 7463
rect 6009 7361 6043 7395
rect 7389 7361 7423 7395
rect 8585 7361 8619 7395
rect 11897 7361 11931 7395
rect 14841 7361 14875 7395
rect 17785 7361 17819 7395
rect 1593 7293 1627 7327
rect 1869 7293 1903 7327
rect 4537 7293 4571 7327
rect 9413 7293 9447 7327
rect 18429 7293 18463 7327
rect 18705 7293 18739 7327
rect 4353 7225 4387 7259
rect 3341 7157 3375 7191
rect 4721 7157 4755 7191
rect 5825 7157 5859 7191
rect 8769 7157 8803 7191
rect 11713 7157 11747 7191
rect 15025 7157 15059 7191
rect 20177 7157 20211 7191
rect 2973 6953 3007 6987
rect 4123 6953 4157 6987
rect 11253 6953 11287 6987
rect 5641 6817 5675 6851
rect 2329 6749 2363 6783
rect 4020 6749 4054 6783
rect 5365 6749 5399 6783
rect 9137 6749 9171 6783
rect 9873 6749 9907 6783
rect 11437 6749 11471 6783
rect 15669 6749 15703 6783
rect 20177 6749 20211 6783
rect 7389 6681 7423 6715
rect 9321 6613 9355 6647
rect 10057 6613 10091 6647
rect 15853 6613 15887 6647
rect 19993 6613 20027 6647
rect 2927 6409 2961 6443
rect 14105 6409 14139 6443
rect 16313 6409 16347 6443
rect 2237 6273 2271 6307
rect 3030 6273 3064 6307
rect 3893 6273 3927 6307
rect 7481 6273 7515 6307
rect 9229 6273 9263 6307
rect 10609 6273 10643 6307
rect 12357 6273 12391 6307
rect 16865 6273 16899 6307
rect 1869 6205 1903 6239
rect 2329 6205 2363 6239
rect 5273 6205 5307 6239
rect 7389 6205 7423 6239
rect 9965 6205 9999 6239
rect 12633 6205 12667 6239
rect 17141 6205 17175 6239
rect 5089 6137 5123 6171
rect 9781 6137 9815 6171
rect 15945 6137 15979 6171
rect 4537 6069 4571 6103
rect 5457 6069 5491 6103
rect 7849 6069 7883 6103
rect 8953 6069 8987 6103
rect 10149 6069 10183 6103
rect 10793 6069 10827 6103
rect 14933 6069 14967 6103
rect 18613 6069 18647 6103
rect 6561 5865 6595 5899
rect 9781 5865 9815 5899
rect 12173 5865 12207 5899
rect 15025 5865 15059 5899
rect 16037 5797 16071 5831
rect 3157 5729 3191 5763
rect 3433 5729 3467 5763
rect 4261 5729 4295 5763
rect 6193 5729 6227 5763
rect 6377 5729 6411 5763
rect 7435 5729 7469 5763
rect 10425 5729 10459 5763
rect 17417 5729 17451 5763
rect 3065 5661 3099 5695
rect 3985 5661 4019 5695
rect 7348 5661 7382 5695
rect 7941 5661 7975 5695
rect 8585 5661 8619 5695
rect 9137 5661 9171 5695
rect 17141 5661 17175 5695
rect 10701 5593 10735 5627
rect 5733 5525 5767 5559
rect 16405 5525 16439 5559
rect 18889 5525 18923 5559
rect 5181 5321 5215 5355
rect 6929 5321 6963 5355
rect 9413 5321 9447 5355
rect 13461 5321 13495 5355
rect 7941 5253 7975 5287
rect 17509 5253 17543 5287
rect 4537 5185 4571 5219
rect 5676 5185 5710 5219
rect 6745 5185 6779 5219
rect 10057 5185 10091 5219
rect 11713 5185 11747 5219
rect 13921 5185 13955 5219
rect 17233 5185 17267 5219
rect 19901 5185 19935 5219
rect 7665 5117 7699 5151
rect 9873 5117 9907 5151
rect 11989 5117 12023 5151
rect 14197 5117 14231 5151
rect 18981 5117 19015 5151
rect 5779 5049 5813 5083
rect 6561 5049 6595 5083
rect 10241 4981 10275 5015
rect 15669 4981 15703 5015
rect 20085 4981 20119 5015
rect 4951 4777 4985 4811
rect 8125 4777 8159 4811
rect 14933 4777 14967 4811
rect 15945 4709 15979 4743
rect 3433 4641 3467 4675
rect 9321 4641 9355 4675
rect 9505 4641 9539 4675
rect 10011 4641 10045 4675
rect 3065 4573 3099 4607
rect 4880 4573 4914 4607
rect 6377 4573 6411 4607
rect 10114 4573 10148 4607
rect 6653 4505 6687 4539
rect 9137 4505 9171 4539
rect 1639 4437 1673 4471
rect 16313 4437 16347 4471
rect 6607 4233 6641 4267
rect 3249 4097 3283 4131
rect 3617 4097 3651 4131
rect 6710 4097 6744 4131
rect 8033 4097 8067 4131
rect 17785 4097 17819 4131
rect 8401 4029 8435 4063
rect 18061 4029 18095 4063
rect 1823 3893 1857 3927
rect 9827 3893 9861 3927
rect 19533 3893 19567 3927
rect 2421 3621 2455 3655
rect 5089 3553 5123 3587
rect 10977 3553 11011 3587
rect 15485 3553 15519 3587
rect 15853 3553 15887 3587
rect 1593 3485 1627 3519
rect 2605 3485 2639 3519
rect 4629 3485 4663 3519
rect 10609 3485 10643 3519
rect 19901 3485 19935 3519
rect 5365 3417 5399 3451
rect 1777 3349 1811 3383
rect 4445 3349 4479 3383
rect 6837 3349 6871 3383
rect 12403 3349 12437 3383
rect 17279 3349 17313 3383
rect 20085 3349 20119 3383
rect 4859 3145 4893 3179
rect 6837 3077 6871 3111
rect 1593 3009 1627 3043
rect 2329 3009 2363 3043
rect 3065 3009 3099 3043
rect 3433 3009 3467 3043
rect 6009 3009 6043 3043
rect 9321 3009 9355 3043
rect 16865 3009 16899 3043
rect 19165 3009 19199 3043
rect 19901 3009 19935 3043
rect 6561 2941 6595 2975
rect 9689 2941 9723 2975
rect 17233 2941 17267 2975
rect 18659 2941 18693 2975
rect 1777 2805 1811 2839
rect 2513 2805 2547 2839
rect 5825 2805 5859 2839
rect 8309 2805 8343 2839
rect 11115 2805 11149 2839
rect 19349 2805 19383 2839
rect 20085 2805 20119 2839
rect 3341 2601 3375 2635
rect 4340 2601 4374 2635
rect 5825 2601 5859 2635
rect 18705 2601 18739 2635
rect 1593 2465 1627 2499
rect 4077 2397 4111 2431
rect 7113 2397 7147 2431
rect 8309 2397 8343 2431
rect 9965 2397 9999 2431
rect 11161 2397 11195 2431
rect 12541 2397 12575 2431
rect 14289 2397 14323 2431
rect 15301 2397 15335 2431
rect 16865 2397 16899 2431
rect 17601 2397 17635 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 1869 2329 1903 2363
rect 7297 2261 7331 2295
rect 8493 2261 8527 2295
rect 9781 2261 9815 2295
rect 10977 2261 11011 2295
rect 12357 2261 12391 2295
rect 14473 2261 14507 2295
rect 15117 2261 15151 2295
rect 17049 2261 17083 2295
rect 17785 2261 17819 2295
rect 19625 2261 19659 2295
<< metal1 >>
rect 1104 21786 20859 21808
rect 1104 21734 5848 21786
rect 5900 21734 5912 21786
rect 5964 21734 5976 21786
rect 6028 21734 6040 21786
rect 6092 21734 6104 21786
rect 6156 21734 10747 21786
rect 10799 21734 10811 21786
rect 10863 21734 10875 21786
rect 10927 21734 10939 21786
rect 10991 21734 11003 21786
rect 11055 21734 15646 21786
rect 15698 21734 15710 21786
rect 15762 21734 15774 21786
rect 15826 21734 15838 21786
rect 15890 21734 15902 21786
rect 15954 21734 20545 21786
rect 20597 21734 20609 21786
rect 20661 21734 20673 21786
rect 20725 21734 20737 21786
rect 20789 21734 20801 21786
rect 20853 21734 20859 21786
rect 1104 21712 20859 21734
rect 1854 21632 1860 21684
rect 1912 21672 1918 21684
rect 2041 21675 2099 21681
rect 2041 21672 2053 21675
rect 1912 21644 2053 21672
rect 1912 21632 1918 21644
rect 2041 21641 2053 21644
rect 2087 21641 2099 21675
rect 2041 21635 2099 21641
rect 3142 21632 3148 21684
rect 3200 21672 3206 21684
rect 3237 21675 3295 21681
rect 3237 21672 3249 21675
rect 3200 21644 3249 21672
rect 3200 21632 3206 21644
rect 3237 21641 3249 21644
rect 3283 21641 3295 21675
rect 4614 21672 4620 21684
rect 4575 21644 4620 21672
rect 3237 21635 3295 21641
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 5905 21675 5963 21681
rect 5905 21672 5917 21675
rect 5776 21644 5917 21672
rect 5776 21632 5782 21644
rect 5905 21641 5917 21644
rect 5951 21641 5963 21675
rect 7282 21672 7288 21684
rect 7243 21644 7288 21672
rect 5905 21635 5963 21641
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 8294 21632 8300 21684
rect 8352 21672 8358 21684
rect 8481 21675 8539 21681
rect 8481 21672 8493 21675
rect 8352 21644 8493 21672
rect 8352 21632 8358 21644
rect 8481 21641 8493 21644
rect 8527 21641 8539 21675
rect 8481 21635 8539 21641
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 9861 21675 9919 21681
rect 9861 21672 9873 21675
rect 9732 21644 9873 21672
rect 9732 21632 9738 21644
rect 9861 21641 9873 21644
rect 9907 21641 9919 21675
rect 9861 21635 9919 21641
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 10965 21675 11023 21681
rect 10965 21672 10977 21675
rect 10652 21644 10977 21672
rect 10652 21632 10658 21644
rect 10965 21641 10977 21644
rect 11011 21641 11023 21675
rect 12342 21672 12348 21684
rect 12303 21644 12348 21672
rect 10965 21635 11023 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 13814 21632 13820 21684
rect 13872 21672 13878 21684
rect 14461 21675 14519 21681
rect 14461 21672 14473 21675
rect 13872 21644 14473 21672
rect 13872 21632 13878 21644
rect 14461 21641 14473 21644
rect 14507 21641 14519 21675
rect 14461 21635 14519 21641
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 15197 21675 15255 21681
rect 15197 21672 15209 21675
rect 14792 21644 15209 21672
rect 14792 21632 14798 21644
rect 15197 21641 15209 21644
rect 15243 21641 15255 21675
rect 15197 21635 15255 21641
rect 16022 21632 16028 21684
rect 16080 21672 16086 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16080 21644 17049 21672
rect 16080 21632 16086 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17037 21635 17095 21641
rect 17310 21632 17316 21684
rect 17368 21672 17374 21684
rect 17773 21675 17831 21681
rect 17773 21672 17785 21675
rect 17368 21644 17785 21672
rect 17368 21632 17374 21644
rect 17773 21641 17785 21644
rect 17819 21641 17831 21675
rect 17773 21635 17831 21641
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 19613 21675 19671 21681
rect 19613 21672 19625 21675
rect 18656 21644 19625 21672
rect 18656 21632 18662 21644
rect 19613 21641 19625 21644
rect 19659 21641 19671 21675
rect 19613 21635 19671 21641
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21536 2283 21539
rect 3234 21536 3240 21548
rect 2271 21508 3240 21536
rect 2271 21505 2283 21508
rect 2225 21499 2283 21505
rect 3234 21496 3240 21508
rect 3292 21496 3298 21548
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21536 3479 21539
rect 4062 21536 4068 21548
rect 3467 21508 4068 21536
rect 3467 21505 3479 21508
rect 3421 21499 3479 21505
rect 4062 21496 4068 21508
rect 4120 21496 4126 21548
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21536 4859 21539
rect 4890 21536 4896 21548
rect 4847 21508 4896 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 5626 21496 5632 21548
rect 5684 21536 5690 21548
rect 5721 21539 5779 21545
rect 5721 21536 5733 21539
rect 5684 21508 5733 21536
rect 5684 21496 5690 21508
rect 5721 21505 5733 21508
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21536 7159 21539
rect 7466 21536 7472 21548
rect 7147 21508 7472 21536
rect 7147 21505 7159 21508
rect 7101 21499 7159 21505
rect 7466 21496 7472 21508
rect 7524 21496 7530 21548
rect 8297 21539 8355 21545
rect 8297 21505 8309 21539
rect 8343 21536 8355 21539
rect 8938 21536 8944 21548
rect 8343 21508 8944 21536
rect 8343 21505 8355 21508
rect 8297 21499 8355 21505
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 9674 21536 9680 21548
rect 9635 21508 9680 21536
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 11146 21536 11152 21548
rect 11107 21508 11152 21536
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 12526 21536 12532 21548
rect 12487 21508 12532 21536
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14277 21539 14335 21545
rect 14277 21536 14289 21539
rect 14240 21508 14289 21536
rect 14240 21496 14246 21508
rect 14277 21505 14289 21508
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 14424 21508 15025 21536
rect 14424 21496 14430 21508
rect 15013 21505 15025 21508
rect 15059 21505 15071 21539
rect 15013 21499 15071 21505
rect 15898 21539 15956 21545
rect 15898 21505 15910 21539
rect 15944 21536 15956 21539
rect 15944 21508 16528 21536
rect 15944 21505 15956 21508
rect 15898 21499 15956 21505
rect 16500 21468 16528 21508
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16632 21508 16865 21536
rect 16632 21496 16638 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 17586 21536 17592 21548
rect 17547 21508 17592 21536
rect 16853 21499 16911 21505
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 18874 21536 18880 21548
rect 18835 21508 18880 21536
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 19116 21508 19441 21536
rect 19116 21496 19122 21508
rect 19429 21505 19441 21508
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 16666 21468 16672 21480
rect 16500 21440 16672 21468
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 18693 21403 18751 21409
rect 18693 21369 18705 21403
rect 18739 21400 18751 21403
rect 21174 21400 21180 21412
rect 18739 21372 21180 21400
rect 18739 21369 18751 21372
rect 18693 21363 18751 21369
rect 21174 21360 21180 21372
rect 21232 21360 21238 21412
rect 15746 21292 15752 21344
rect 15804 21341 15810 21344
rect 15804 21335 15853 21341
rect 15804 21301 15807 21335
rect 15841 21301 15853 21335
rect 15804 21295 15853 21301
rect 15804 21292 15810 21295
rect 1104 21242 20700 21264
rect 1104 21190 3399 21242
rect 3451 21190 3463 21242
rect 3515 21190 3527 21242
rect 3579 21190 3591 21242
rect 3643 21190 3655 21242
rect 3707 21190 8298 21242
rect 8350 21190 8362 21242
rect 8414 21190 8426 21242
rect 8478 21190 8490 21242
rect 8542 21190 8554 21242
rect 8606 21190 13197 21242
rect 13249 21190 13261 21242
rect 13313 21190 13325 21242
rect 13377 21190 13389 21242
rect 13441 21190 13453 21242
rect 13505 21190 18096 21242
rect 18148 21190 18160 21242
rect 18212 21190 18224 21242
rect 18276 21190 18288 21242
rect 18340 21190 18352 21242
rect 18404 21190 20700 21242
rect 1104 21168 20700 21190
rect 566 21088 572 21140
rect 624 21128 630 21140
rect 1765 21131 1823 21137
rect 1765 21128 1777 21131
rect 624 21100 1777 21128
rect 624 21088 630 21100
rect 1765 21097 1777 21100
rect 1811 21097 1823 21131
rect 14274 21128 14280 21140
rect 1765 21091 1823 21097
rect 6886 21100 14280 21128
rect 6273 20995 6331 21001
rect 6273 20961 6285 20995
rect 6319 20992 6331 20995
rect 6886 20992 6914 21100
rect 14274 21088 14280 21100
rect 14332 21088 14338 21140
rect 17175 21131 17233 21137
rect 17175 21097 17187 21131
rect 17221 21128 17233 21131
rect 17586 21128 17592 21140
rect 17221 21100 17592 21128
rect 17221 21097 17233 21100
rect 17175 21091 17233 21097
rect 17586 21088 17592 21100
rect 17644 21088 17650 21140
rect 19886 21088 19892 21140
rect 19944 21128 19950 21140
rect 20073 21131 20131 21137
rect 20073 21128 20085 21131
rect 19944 21100 20085 21128
rect 19944 21088 19950 21100
rect 20073 21097 20085 21100
rect 20119 21097 20131 21131
rect 20073 21091 20131 21097
rect 13725 20995 13783 21001
rect 13725 20992 13737 20995
rect 6319 20964 6914 20992
rect 7208 20964 13737 20992
rect 6319 20961 6331 20964
rect 6273 20955 6331 20961
rect 1578 20924 1584 20936
rect 1539 20896 1584 20924
rect 1578 20884 1584 20896
rect 1636 20884 1642 20936
rect 2682 20924 2688 20936
rect 2643 20896 2688 20924
rect 2682 20884 2688 20896
rect 2740 20884 2746 20936
rect 6546 20884 6552 20936
rect 6604 20924 6610 20936
rect 7208 20933 7236 20964
rect 13725 20961 13737 20964
rect 13771 20992 13783 20995
rect 15746 20992 15752 21004
rect 13771 20964 15608 20992
rect 15707 20964 15752 20992
rect 13771 20961 13783 20964
rect 13725 20955 13783 20961
rect 7009 20927 7067 20933
rect 7009 20924 7021 20927
rect 6604 20896 7021 20924
rect 6604 20884 6610 20896
rect 7009 20893 7021 20896
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20893 7251 20927
rect 7193 20887 7251 20893
rect 8180 20927 8238 20933
rect 8180 20893 8192 20927
rect 8226 20924 8238 20927
rect 9490 20924 9496 20936
rect 8226 20896 9496 20924
rect 8226 20893 8238 20896
rect 8180 20887 8238 20893
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 10134 20924 10140 20936
rect 10095 20896 10140 20924
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 13446 20924 13452 20936
rect 13407 20896 13452 20924
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 15286 20884 15292 20936
rect 15344 20924 15350 20936
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 15344 20896 15393 20924
rect 15344 20884 15350 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15580 20924 15608 20964
rect 15746 20952 15752 20964
rect 15804 20952 15810 21004
rect 19242 20992 19248 21004
rect 15856 20964 19248 20992
rect 15856 20924 15884 20964
rect 19242 20952 19248 20964
rect 19300 20952 19306 21004
rect 15580 20896 15884 20924
rect 15381 20887 15439 20893
rect 16666 20884 16672 20936
rect 16724 20924 16730 20936
rect 17830 20927 17888 20933
rect 17830 20924 17842 20927
rect 16724 20896 17842 20924
rect 16724 20884 16730 20896
rect 17830 20893 17842 20896
rect 17876 20924 17888 20927
rect 18414 20924 18420 20936
rect 18472 20933 18478 20936
rect 18472 20927 18500 20933
rect 17876 20896 18420 20924
rect 17876 20893 17888 20896
rect 17830 20887 17888 20893
rect 18414 20884 18420 20896
rect 18488 20893 18500 20927
rect 19886 20924 19892 20936
rect 19847 20896 19892 20924
rect 18472 20887 18500 20893
rect 18472 20884 18478 20887
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 2774 20816 2780 20868
rect 2832 20856 2838 20868
rect 3237 20859 3295 20865
rect 3237 20856 3249 20859
rect 2832 20828 3249 20856
rect 2832 20816 2838 20828
rect 3237 20825 3249 20828
rect 3283 20856 3295 20859
rect 3878 20856 3884 20868
rect 3283 20828 3884 20856
rect 3283 20825 3295 20828
rect 3237 20819 3295 20825
rect 3878 20816 3884 20828
rect 3936 20816 3942 20868
rect 6914 20856 6920 20868
rect 5842 20828 6920 20856
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 10410 20856 10416 20868
rect 10371 20828 10416 20856
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 11422 20816 11428 20868
rect 11480 20816 11486 20868
rect 17586 20856 17592 20868
rect 16790 20828 17592 20856
rect 17586 20816 17592 20828
rect 17644 20816 17650 20868
rect 4801 20791 4859 20797
rect 4801 20757 4813 20791
rect 4847 20788 4859 20791
rect 5534 20788 5540 20800
rect 4847 20760 5540 20788
rect 4847 20757 4859 20760
rect 4801 20751 4859 20757
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 8294 20797 8300 20800
rect 8251 20791 8300 20797
rect 8251 20757 8263 20791
rect 8297 20757 8300 20791
rect 8251 20751 8300 20757
rect 8294 20748 8300 20751
rect 8352 20748 8358 20800
rect 11330 20748 11336 20800
rect 11388 20788 11394 20800
rect 11885 20791 11943 20797
rect 11885 20788 11897 20791
rect 11388 20760 11897 20788
rect 11388 20748 11394 20760
rect 11885 20757 11897 20760
rect 11931 20757 11943 20791
rect 11885 20751 11943 20757
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17727 20791 17785 20797
rect 17727 20788 17739 20791
rect 17276 20760 17739 20788
rect 17276 20748 17282 20760
rect 17727 20757 17739 20760
rect 17773 20757 17785 20791
rect 17727 20751 17785 20757
rect 17862 20748 17868 20800
rect 17920 20788 17926 20800
rect 18371 20791 18429 20797
rect 18371 20788 18383 20791
rect 17920 20760 18383 20788
rect 17920 20748 17926 20760
rect 18371 20757 18383 20760
rect 18417 20757 18429 20791
rect 18371 20751 18429 20757
rect 1104 20698 20859 20720
rect 1104 20646 5848 20698
rect 5900 20646 5912 20698
rect 5964 20646 5976 20698
rect 6028 20646 6040 20698
rect 6092 20646 6104 20698
rect 6156 20646 10747 20698
rect 10799 20646 10811 20698
rect 10863 20646 10875 20698
rect 10927 20646 10939 20698
rect 10991 20646 11003 20698
rect 11055 20646 15646 20698
rect 15698 20646 15710 20698
rect 15762 20646 15774 20698
rect 15826 20646 15838 20698
rect 15890 20646 15902 20698
rect 15954 20646 20545 20698
rect 20597 20646 20609 20698
rect 20661 20646 20673 20698
rect 20725 20646 20737 20698
rect 20789 20646 20801 20698
rect 20853 20646 20859 20698
rect 1104 20624 20859 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 9674 20544 9680 20596
rect 9732 20593 9738 20596
rect 9732 20587 9781 20593
rect 9732 20553 9735 20587
rect 9769 20553 9781 20587
rect 13446 20584 13452 20596
rect 9732 20547 9781 20553
rect 11900 20556 13452 20584
rect 9732 20544 9738 20547
rect 2774 20516 2780 20528
rect 1872 20488 2780 20516
rect 1872 20457 1900 20488
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 4246 20476 4252 20528
rect 4304 20476 4310 20528
rect 4709 20519 4767 20525
rect 4709 20485 4721 20519
rect 4755 20516 4767 20519
rect 5859 20519 5917 20525
rect 5859 20516 5871 20519
rect 4755 20488 5871 20516
rect 4755 20485 4767 20488
rect 4709 20479 4767 20485
rect 5859 20485 5871 20488
rect 5905 20485 5917 20519
rect 9858 20516 9864 20528
rect 9338 20488 9864 20516
rect 5859 20479 5917 20485
rect 9858 20476 9864 20488
rect 9916 20476 9922 20528
rect 11900 20516 11928 20556
rect 13446 20544 13452 20556
rect 13504 20544 13510 20596
rect 13541 20587 13599 20593
rect 13541 20553 13553 20587
rect 13587 20584 13599 20587
rect 18647 20587 18705 20593
rect 13587 20556 14320 20584
rect 13587 20553 13599 20556
rect 13541 20547 13599 20553
rect 14292 20525 14320 20556
rect 18647 20553 18659 20587
rect 18693 20584 18705 20587
rect 19058 20584 19064 20596
rect 18693 20556 19064 20584
rect 18693 20553 18705 20556
rect 18647 20547 18705 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19242 20584 19248 20596
rect 19203 20556 19248 20584
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 11808 20488 11928 20516
rect 14277 20519 14335 20525
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20417 1915 20451
rect 2590 20448 2596 20460
rect 2551 20420 2596 20448
rect 1857 20411 1915 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 5962 20451 6020 20457
rect 5962 20417 5974 20451
rect 6008 20448 6020 20451
rect 7282 20448 7288 20460
rect 6008 20420 7288 20448
rect 6008 20417 6020 20420
rect 5962 20411 6020 20417
rect 7282 20408 7288 20420
rect 7340 20408 7346 20460
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20448 7435 20451
rect 8018 20448 8024 20460
rect 7423 20420 8024 20448
rect 7423 20417 7435 20420
rect 7377 20411 7435 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8294 20448 8300 20460
rect 8255 20420 8300 20448
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 10134 20408 10140 20460
rect 10192 20448 10198 20460
rect 11054 20448 11060 20460
rect 10192 20420 11060 20448
rect 10192 20408 10198 20420
rect 11054 20408 11060 20420
rect 11112 20448 11118 20460
rect 11808 20457 11836 20488
rect 14277 20485 14289 20519
rect 14323 20485 14335 20519
rect 14277 20479 14335 20485
rect 17586 20476 17592 20528
rect 17644 20476 17650 20528
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11112 20420 11805 20448
rect 11112 20408 11118 20420
rect 11793 20417 11805 20420
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 2608 20380 2636 20408
rect 3237 20383 3295 20389
rect 3237 20380 3249 20383
rect 2608 20352 3249 20380
rect 3237 20349 3249 20352
rect 3283 20349 3295 20383
rect 3237 20343 3295 20349
rect 4985 20383 5043 20389
rect 4985 20349 4997 20383
rect 5031 20380 5043 20383
rect 5718 20380 5724 20392
rect 5031 20352 5724 20380
rect 5031 20349 5043 20352
rect 4985 20343 5043 20349
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20380 7987 20383
rect 10318 20380 10324 20392
rect 7975 20352 10324 20380
rect 7975 20349 7987 20352
rect 7929 20343 7987 20349
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20380 12127 20383
rect 12802 20380 12808 20392
rect 12115 20352 12808 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 2774 20244 2780 20256
rect 2735 20216 2780 20244
rect 2774 20204 2780 20216
rect 2832 20204 2838 20256
rect 4246 20204 4252 20256
rect 4304 20244 4310 20256
rect 7006 20244 7012 20256
rect 4304 20216 7012 20244
rect 4304 20204 4310 20216
rect 7006 20204 7012 20216
rect 7064 20244 7070 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 7064 20216 7113 20244
rect 7064 20204 7070 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 13188 20244 13216 20434
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 19426 20448 19432 20460
rect 19387 20420 19432 20448
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 19576 20420 19901 20448
rect 19576 20408 19582 20420
rect 19889 20417 19901 20420
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14001 20383 14059 20389
rect 14001 20380 14013 20383
rect 13504 20352 14013 20380
rect 13504 20340 13510 20352
rect 14001 20349 14013 20352
rect 14047 20380 14059 20383
rect 16022 20380 16028 20392
rect 14047 20352 16028 20380
rect 14047 20349 14059 20352
rect 14001 20343 14059 20349
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 16758 20340 16764 20392
rect 16816 20380 16822 20392
rect 16853 20383 16911 20389
rect 16853 20380 16865 20383
rect 16816 20352 16865 20380
rect 16816 20340 16822 20352
rect 16853 20349 16865 20352
rect 16899 20349 16911 20383
rect 16853 20343 16911 20349
rect 15470 20244 15476 20256
rect 12492 20216 15476 20244
rect 12492 20204 12498 20216
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 15746 20244 15752 20256
rect 15707 20216 15752 20244
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 20070 20244 20076 20256
rect 20031 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 1104 20154 20700 20176
rect 1104 20102 3399 20154
rect 3451 20102 3463 20154
rect 3515 20102 3527 20154
rect 3579 20102 3591 20154
rect 3643 20102 3655 20154
rect 3707 20102 8298 20154
rect 8350 20102 8362 20154
rect 8414 20102 8426 20154
rect 8478 20102 8490 20154
rect 8542 20102 8554 20154
rect 8606 20102 13197 20154
rect 13249 20102 13261 20154
rect 13313 20102 13325 20154
rect 13377 20102 13389 20154
rect 13441 20102 13453 20154
rect 13505 20102 18096 20154
rect 18148 20102 18160 20154
rect 18212 20102 18224 20154
rect 18276 20102 18288 20154
rect 18340 20102 18352 20154
rect 18404 20102 20700 20154
rect 1104 20080 20700 20102
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 2682 20040 2688 20052
rect 2639 20012 2688 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 2682 20000 2688 20012
rect 2740 20000 2746 20052
rect 7282 20000 7288 20052
rect 7340 20040 7346 20052
rect 7745 20043 7803 20049
rect 7745 20040 7757 20043
rect 7340 20012 7757 20040
rect 7340 20000 7346 20012
rect 7745 20009 7757 20012
rect 7791 20009 7803 20043
rect 12802 20040 12808 20052
rect 12763 20012 12808 20040
rect 7745 20003 7803 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 14274 20040 14280 20052
rect 14235 20012 14280 20040
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 5592 19876 6285 19904
rect 5592 19864 5598 19876
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6273 19867 6331 19873
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 11054 19904 11060 19916
rect 9272 19876 11060 19904
rect 9272 19864 9278 19876
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11330 19904 11336 19916
rect 11291 19876 11336 19904
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 15746 19904 15752 19916
rect 15707 19876 15752 19904
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 16022 19904 16028 19916
rect 15983 19876 16028 19904
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 17405 19907 17463 19913
rect 17405 19873 17417 19907
rect 17451 19904 17463 19907
rect 17862 19904 17868 19916
rect 17451 19876 17868 19904
rect 17451 19873 17463 19876
rect 17405 19867 17463 19873
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 2774 19836 2780 19848
rect 2735 19808 2780 19836
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 5997 19839 6055 19845
rect 5997 19836 6009 19839
rect 5776 19808 6009 19836
rect 5776 19796 5782 19808
rect 5997 19805 6009 19808
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 6012 19768 6040 19799
rect 12434 19796 12440 19848
rect 12492 19796 12498 19848
rect 16482 19836 16488 19848
rect 16443 19808 16488 19836
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 17126 19836 17132 19848
rect 17087 19808 17132 19836
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 18932 19808 19625 19836
rect 18932 19796 18938 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 6546 19768 6552 19780
rect 6012 19740 6552 19768
rect 6546 19728 6552 19740
rect 6604 19728 6610 19780
rect 7006 19728 7012 19780
rect 7064 19728 7070 19780
rect 15470 19768 15476 19780
rect 15318 19740 15476 19768
rect 15470 19728 15476 19740
rect 15528 19768 15534 19780
rect 17034 19768 17040 19780
rect 15528 19740 17040 19768
rect 15528 19728 15534 19740
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 18966 19768 18972 19780
rect 18630 19740 18972 19768
rect 18966 19728 18972 19740
rect 19024 19768 19030 19780
rect 19797 19771 19855 19777
rect 19797 19768 19809 19771
rect 19024 19740 19809 19768
rect 19024 19728 19030 19740
rect 19797 19737 19809 19740
rect 19843 19737 19855 19771
rect 19797 19731 19855 19737
rect 8018 19660 8024 19712
rect 8076 19700 8082 19712
rect 11238 19700 11244 19712
rect 8076 19672 11244 19700
rect 8076 19660 8082 19672
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19700 16727 19703
rect 18690 19700 18696 19712
rect 16715 19672 18696 19700
rect 16715 19669 16727 19672
rect 16669 19663 16727 19669
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 1104 19610 20859 19632
rect 1104 19558 5848 19610
rect 5900 19558 5912 19610
rect 5964 19558 5976 19610
rect 6028 19558 6040 19610
rect 6092 19558 6104 19610
rect 6156 19558 10747 19610
rect 10799 19558 10811 19610
rect 10863 19558 10875 19610
rect 10927 19558 10939 19610
rect 10991 19558 11003 19610
rect 11055 19558 15646 19610
rect 15698 19558 15710 19610
rect 15762 19558 15774 19610
rect 15826 19558 15838 19610
rect 15890 19558 15902 19610
rect 15954 19558 20545 19610
rect 20597 19558 20609 19610
rect 20661 19558 20673 19610
rect 20725 19558 20737 19610
rect 20789 19558 20801 19610
rect 20853 19558 20859 19610
rect 1104 19536 20859 19558
rect 7009 19499 7067 19505
rect 7009 19465 7021 19499
rect 7055 19496 7067 19499
rect 7055 19468 9536 19496
rect 7055 19465 7067 19468
rect 7009 19459 7067 19465
rect 2590 19428 2596 19440
rect 2551 19400 2596 19428
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 4246 19428 4252 19440
rect 3818 19400 4252 19428
rect 4246 19388 4252 19400
rect 4304 19388 4310 19440
rect 8018 19388 8024 19440
rect 8076 19388 8082 19440
rect 9508 19437 9536 19468
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10468 19468 10977 19496
rect 10468 19456 10474 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 17635 19499 17693 19505
rect 17635 19465 17647 19499
rect 17681 19496 17693 19499
rect 19426 19496 19432 19508
rect 17681 19468 19432 19496
rect 17681 19465 17693 19468
rect 17635 19459 17693 19465
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 9493 19431 9551 19437
rect 9493 19397 9505 19431
rect 9539 19397 9551 19431
rect 11238 19428 11244 19440
rect 10718 19400 11244 19428
rect 9493 19391 9551 19397
rect 11238 19388 11244 19400
rect 11296 19388 11302 19440
rect 18966 19388 18972 19440
rect 19024 19388 19030 19440
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19360 8815 19363
rect 9214 19360 9220 19372
rect 8803 19332 9220 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16888 19363 16946 19369
rect 16888 19360 16900 19363
rect 16264 19332 16900 19360
rect 16264 19320 16270 19332
rect 16888 19329 16900 19332
rect 16934 19329 16946 19363
rect 16888 19323 16946 19329
rect 17564 19363 17622 19369
rect 17564 19329 17576 19363
rect 17610 19360 17622 19363
rect 17862 19360 17868 19372
rect 17610 19332 17868 19360
rect 17610 19329 17622 19332
rect 17564 19323 17622 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 8481 19295 8539 19301
rect 8481 19261 8493 19295
rect 8527 19292 8539 19295
rect 8527 19264 8708 19292
rect 8527 19261 8539 19264
rect 8481 19255 8539 19261
rect 8680 19168 8708 19264
rect 17126 19252 17132 19304
rect 17184 19292 17190 19304
rect 17954 19292 17960 19304
rect 17184 19264 17960 19292
rect 17184 19252 17190 19264
rect 17954 19252 17960 19264
rect 18012 19292 18018 19304
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 18012 19264 18245 19292
rect 18012 19252 18018 19264
rect 18233 19261 18245 19264
rect 18279 19261 18291 19295
rect 18506 19292 18512 19304
rect 18467 19264 18512 19292
rect 18233 19255 18291 19261
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 4065 19159 4123 19165
rect 4065 19125 4077 19159
rect 4111 19156 4123 19159
rect 4246 19156 4252 19168
rect 4111 19128 4252 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 16991 19159 17049 19165
rect 16991 19125 17003 19159
rect 17037 19156 17049 19159
rect 17218 19156 17224 19168
rect 17037 19128 17224 19156
rect 17037 19125 17049 19128
rect 16991 19119 17049 19125
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 19702 19116 19708 19168
rect 19760 19156 19766 19168
rect 19981 19159 20039 19165
rect 19981 19156 19993 19159
rect 19760 19128 19993 19156
rect 19760 19116 19766 19128
rect 19981 19125 19993 19128
rect 20027 19125 20039 19159
rect 19981 19119 20039 19125
rect 1104 19066 20700 19088
rect 1104 19014 3399 19066
rect 3451 19014 3463 19066
rect 3515 19014 3527 19066
rect 3579 19014 3591 19066
rect 3643 19014 3655 19066
rect 3707 19014 8298 19066
rect 8350 19014 8362 19066
rect 8414 19014 8426 19066
rect 8478 19014 8490 19066
rect 8542 19014 8554 19066
rect 8606 19014 13197 19066
rect 13249 19014 13261 19066
rect 13313 19014 13325 19066
rect 13377 19014 13389 19066
rect 13441 19014 13453 19066
rect 13505 19014 18096 19066
rect 18148 19014 18160 19066
rect 18212 19014 18224 19066
rect 18276 19014 18288 19066
rect 18340 19014 18352 19066
rect 18404 19014 20700 19066
rect 1104 18992 20700 19014
rect 8573 18955 8631 18961
rect 8573 18921 8585 18955
rect 8619 18952 8631 18955
rect 8662 18952 8668 18964
rect 8619 18924 8668 18952
rect 8619 18921 8631 18924
rect 8573 18915 8631 18921
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 12526 18961 12532 18964
rect 12483 18955 12532 18961
rect 12483 18921 12495 18955
rect 12529 18921 12532 18955
rect 12483 18915 12532 18921
rect 12526 18912 12532 18915
rect 12584 18912 12590 18964
rect 17862 18952 17868 18964
rect 17823 18924 17868 18952
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 17034 18844 17040 18896
rect 17092 18884 17098 18896
rect 19794 18884 19800 18896
rect 17092 18856 19800 18884
rect 17092 18844 17098 18856
rect 19794 18844 19800 18856
rect 19852 18844 19858 18896
rect 2314 18776 2320 18828
rect 2372 18816 2378 18828
rect 3973 18819 4031 18825
rect 3973 18816 3985 18819
rect 2372 18788 3985 18816
rect 2372 18776 2378 18788
rect 3973 18785 3985 18788
rect 4019 18785 4031 18819
rect 4246 18816 4252 18828
rect 4207 18788 4252 18816
rect 3973 18779 4031 18785
rect 3988 18612 4016 18779
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 11057 18819 11115 18825
rect 11057 18785 11069 18819
rect 11103 18816 11115 18819
rect 12434 18816 12440 18828
rect 11103 18788 12440 18816
rect 11103 18785 11115 18788
rect 11057 18779 11115 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 16206 18776 16212 18828
rect 16264 18816 16270 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16264 18788 17509 18816
rect 16264 18776 16270 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 6825 18751 6883 18757
rect 6825 18748 6837 18751
rect 6604 18720 6837 18748
rect 6604 18708 6610 18720
rect 6825 18717 6837 18720
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15378 18748 15384 18760
rect 15335 18720 15384 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 7098 18680 7104 18692
rect 4396 18652 4738 18680
rect 7059 18652 7104 18680
rect 4396 18640 4402 18652
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 7558 18680 7564 18692
rect 7208 18652 7564 18680
rect 5074 18612 5080 18624
rect 3988 18584 5080 18612
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 5721 18615 5779 18621
rect 5721 18612 5733 18615
rect 5684 18584 5733 18612
rect 5684 18572 5690 18584
rect 5721 18581 5733 18584
rect 5767 18581 5779 18615
rect 5721 18575 5779 18581
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 7208 18612 7236 18652
rect 7558 18640 7564 18652
rect 7616 18640 7622 18692
rect 7064 18584 7236 18612
rect 10704 18612 10732 18711
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15979 18720 16405 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 17034 18748 17040 18760
rect 16947 18720 17040 18748
rect 16393 18711 16451 18717
rect 17034 18708 17040 18720
rect 17092 18748 17098 18760
rect 18506 18757 18512 18760
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17092 18720 17693 18748
rect 17092 18708 17098 18720
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 18474 18751 18512 18757
rect 18474 18717 18486 18751
rect 18474 18711 18512 18717
rect 18506 18708 18512 18711
rect 18564 18708 18570 18760
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18748 20223 18751
rect 20254 18748 20260 18760
rect 20211 18720 20260 18748
rect 20211 18717 20223 18720
rect 20165 18711 20223 18717
rect 20254 18708 20260 18720
rect 20312 18708 20318 18760
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 16022 18680 16028 18692
rect 12124 18652 16028 18680
rect 12124 18640 12130 18652
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 11698 18612 11704 18624
rect 10704 18584 11704 18612
rect 7064 18572 7070 18584
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 18371 18615 18429 18621
rect 18371 18612 18383 18615
rect 18196 18584 18383 18612
rect 18196 18572 18202 18584
rect 18371 18581 18383 18584
rect 18417 18581 18429 18615
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 18371 18575 18429 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 1104 18540 20859 18544
rect 1104 18460 1120 18540
rect 1470 18522 20859 18540
rect 1470 18470 5848 18522
rect 5900 18470 5912 18522
rect 5964 18470 5976 18522
rect 6028 18470 6040 18522
rect 6092 18470 6104 18522
rect 6156 18470 10747 18522
rect 10799 18470 10811 18522
rect 10863 18470 10875 18522
rect 10927 18470 10939 18522
rect 10991 18470 11003 18522
rect 11055 18470 15646 18522
rect 15698 18470 15710 18522
rect 15762 18470 15774 18522
rect 15826 18470 15838 18522
rect 15890 18470 15902 18522
rect 15954 18470 20545 18522
rect 20597 18470 20609 18522
rect 20661 18470 20673 18522
rect 20725 18470 20737 18522
rect 20789 18470 20801 18522
rect 20853 18470 20859 18522
rect 1470 18460 20859 18470
rect 1104 18448 20859 18460
rect 7006 18408 7012 18420
rect 4540 18380 7012 18408
rect 4540 18284 4568 18380
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 7098 18368 7104 18420
rect 7156 18408 7162 18420
rect 11146 18417 11152 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 7156 18380 8309 18408
rect 7156 18368 7162 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 11103 18411 11152 18417
rect 11103 18377 11115 18411
rect 11149 18377 11152 18411
rect 11103 18371 11152 18377
rect 11146 18368 11152 18371
rect 11204 18368 11210 18420
rect 12434 18368 12440 18420
rect 12492 18417 12498 18420
rect 12492 18411 12541 18417
rect 12492 18377 12495 18411
rect 12529 18377 12541 18411
rect 15378 18408 15384 18420
rect 12492 18371 12541 18377
rect 14476 18380 15384 18408
rect 12492 18368 12498 18371
rect 5626 18340 5632 18352
rect 5587 18312 5632 18340
rect 5626 18300 5632 18312
rect 5684 18300 5690 18352
rect 7558 18300 7564 18352
rect 7616 18300 7622 18352
rect 12066 18340 12072 18352
rect 10718 18312 12072 18340
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 2501 18275 2559 18281
rect 2501 18272 2513 18275
rect 2372 18244 2513 18272
rect 2372 18232 2378 18244
rect 2501 18241 2513 18244
rect 2547 18241 2559 18275
rect 2501 18235 2559 18241
rect 4522 18232 4528 18284
rect 4580 18232 4586 18284
rect 9309 18275 9367 18281
rect 9309 18241 9321 18275
rect 9355 18272 9367 18275
rect 11977 18275 12035 18281
rect 9355 18244 9812 18272
rect 9355 18241 9367 18244
rect 9309 18235 9367 18241
rect 5074 18164 5080 18216
rect 5132 18204 5138 18216
rect 5905 18207 5963 18213
rect 5905 18204 5917 18207
rect 5132 18176 5917 18204
rect 5132 18164 5138 18176
rect 5905 18173 5917 18176
rect 5951 18204 5963 18207
rect 6546 18204 6552 18216
rect 5951 18176 6552 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 6546 18164 6552 18176
rect 6604 18164 6610 18216
rect 6822 18204 6828 18216
rect 6783 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 9674 18204 9680 18216
rect 9635 18176 9680 18204
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 9784 18204 9812 18244
rect 11977 18241 11989 18275
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 10226 18204 10232 18216
rect 9784 18176 10232 18204
rect 10226 18164 10232 18176
rect 10284 18164 10290 18216
rect 11992 18204 12020 18235
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 14476 18281 14504 18380
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 16206 18408 16212 18420
rect 16167 18380 16212 18408
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 18874 18408 18880 18420
rect 16408 18380 18880 18408
rect 16022 18340 16028 18352
rect 15935 18312 16028 18340
rect 16022 18300 16028 18312
rect 16080 18340 16086 18352
rect 16408 18340 16436 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 19886 18408 19892 18420
rect 19659 18380 19892 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 19886 18368 19892 18380
rect 19944 18368 19950 18420
rect 18138 18340 18144 18352
rect 16080 18312 16436 18340
rect 18099 18312 18144 18340
rect 16080 18300 16086 18312
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 18782 18300 18788 18352
rect 18840 18300 18846 18352
rect 12554 18275 12612 18281
rect 12554 18272 12566 18275
rect 12492 18244 12566 18272
rect 12492 18232 12498 18244
rect 12554 18241 12566 18244
rect 12600 18241 12612 18275
rect 12554 18235 12612 18241
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 17034 18272 17040 18284
rect 16995 18244 17040 18272
rect 14461 18235 14519 18241
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 14274 18204 14280 18216
rect 11992 18176 14280 18204
rect 14274 18164 14280 18176
rect 14332 18164 14338 18216
rect 14734 18204 14740 18216
rect 14695 18176 14740 18204
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 17218 18204 17224 18216
rect 17179 18176 17224 18204
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 17862 18204 17868 18216
rect 17823 18176 17868 18204
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 1857 18071 1915 18077
rect 1857 18037 1869 18071
rect 1903 18068 1915 18071
rect 1946 18068 1952 18080
rect 1903 18040 1952 18068
rect 1903 18037 1915 18040
rect 1857 18031 1915 18037
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 4154 18068 4160 18080
rect 4115 18040 4160 18068
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 11793 18071 11851 18077
rect 11793 18037 11805 18071
rect 11839 18068 11851 18071
rect 12434 18068 12440 18080
rect 11839 18040 12440 18068
rect 11839 18037 11851 18040
rect 11793 18031 11851 18037
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16816 18040 16865 18068
rect 16816 18028 16822 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 1104 17978 20700 18000
rect 1104 17926 3399 17978
rect 3451 17926 3463 17978
rect 3515 17926 3527 17978
rect 3579 17926 3591 17978
rect 3643 17926 3655 17978
rect 3707 17926 8298 17978
rect 8350 17926 8362 17978
rect 8414 17926 8426 17978
rect 8478 17926 8490 17978
rect 8542 17926 8554 17978
rect 8606 17926 13197 17978
rect 13249 17926 13261 17978
rect 13313 17926 13325 17978
rect 13377 17926 13389 17978
rect 13441 17926 13453 17978
rect 13505 17926 18096 17978
rect 18148 17926 18160 17978
rect 18212 17926 18224 17978
rect 18276 17926 18288 17978
rect 18340 17926 18352 17978
rect 18404 17926 20700 17978
rect 1104 17904 20700 17926
rect 6822 17864 6828 17876
rect 6783 17836 6828 17864
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 9674 17873 9680 17876
rect 9631 17867 9680 17873
rect 9631 17833 9643 17867
rect 9677 17833 9680 17867
rect 9631 17827 9680 17833
rect 9674 17824 9680 17827
rect 9732 17824 9738 17876
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 11296 17836 14688 17864
rect 11296 17824 11302 17836
rect 14660 17796 14688 17836
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 14829 17867 14887 17873
rect 14829 17864 14841 17867
rect 14792 17836 14841 17864
rect 14792 17824 14798 17836
rect 14829 17833 14841 17836
rect 14875 17833 14887 17867
rect 14829 17827 14887 17833
rect 17083 17867 17141 17873
rect 17083 17833 17095 17867
rect 17129 17864 17141 17867
rect 19518 17864 19524 17876
rect 17129 17836 19524 17864
rect 17129 17833 17141 17836
rect 17083 17827 17141 17833
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 14660 17768 18920 17796
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 5353 17731 5411 17737
rect 5353 17728 5365 17731
rect 4212 17700 5365 17728
rect 4212 17688 4218 17700
rect 5353 17697 5365 17700
rect 5399 17697 5411 17731
rect 5353 17691 5411 17697
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17728 12035 17731
rect 12434 17728 12440 17740
rect 12023 17700 12440 17728
rect 12023 17697 12035 17700
rect 11977 17691 12035 17697
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 14090 17688 14096 17740
rect 14148 17728 14154 17740
rect 14274 17728 14280 17740
rect 14148 17700 14280 17728
rect 14148 17688 14154 17700
rect 14274 17688 14280 17700
rect 14332 17728 14338 17740
rect 14369 17731 14427 17737
rect 14369 17728 14381 17731
rect 14332 17700 14381 17728
rect 14332 17688 14338 17700
rect 14369 17697 14381 17700
rect 14415 17697 14427 17731
rect 17586 17728 17592 17740
rect 17547 17700 17592 17728
rect 14369 17691 14427 17697
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 17770 17728 17776 17740
rect 17731 17700 17776 17728
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 1946 17660 1952 17672
rect 1907 17632 1952 17660
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2682 17620 2688 17672
rect 2740 17660 2746 17672
rect 3202 17663 3260 17669
rect 3202 17660 3214 17663
rect 2740 17632 3214 17660
rect 2740 17620 2746 17632
rect 3202 17629 3214 17632
rect 3248 17660 3260 17663
rect 5074 17660 5080 17672
rect 3248 17632 4200 17660
rect 5035 17632 5080 17660
rect 3248 17629 3260 17632
rect 3202 17623 3260 17629
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 2593 17527 2651 17533
rect 2593 17524 2605 17527
rect 2556 17496 2605 17524
rect 2556 17484 2562 17496
rect 2593 17493 2605 17496
rect 2639 17493 2651 17527
rect 2593 17487 2651 17493
rect 3050 17484 3056 17536
rect 3108 17533 3114 17536
rect 3108 17527 3157 17533
rect 3108 17493 3111 17527
rect 3145 17493 3157 17527
rect 4172 17524 4200 17632
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 9490 17660 9496 17672
rect 9548 17669 9554 17672
rect 9548 17663 9586 17669
rect 6886 17632 9496 17660
rect 4522 17552 4528 17604
rect 4580 17592 4586 17604
rect 4580 17564 5842 17592
rect 4580 17552 4586 17564
rect 6886 17524 6914 17632
rect 9490 17620 9496 17632
rect 9574 17629 9586 17663
rect 9548 17623 9586 17629
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17629 11759 17663
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 11701 17623 11759 17629
rect 9548 17620 9554 17623
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 10505 17595 10563 17601
rect 10505 17592 10517 17595
rect 9732 17564 10517 17592
rect 9732 17552 9738 17564
rect 10505 17561 10517 17564
rect 10551 17561 10563 17595
rect 10505 17555 10563 17561
rect 10689 17595 10747 17601
rect 10689 17561 10701 17595
rect 10735 17592 10747 17595
rect 11716 17592 11744 17623
rect 13722 17620 13728 17632
rect 13780 17660 13786 17672
rect 14461 17663 14519 17669
rect 14461 17660 14473 17663
rect 13780 17632 14473 17660
rect 13780 17620 13786 17632
rect 14461 17629 14473 17632
rect 14507 17629 14519 17663
rect 14461 17623 14519 17629
rect 17012 17663 17070 17669
rect 17012 17629 17024 17663
rect 17058 17660 17070 17663
rect 17678 17660 17684 17672
rect 17058 17632 17684 17660
rect 17058 17629 17070 17632
rect 17012 17623 17070 17629
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 18690 17660 18696 17672
rect 18651 17632 18696 17660
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 18892 17669 18920 17768
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17660 18935 17663
rect 18923 17632 20116 17660
rect 18923 17629 18935 17632
rect 18877 17623 18935 17629
rect 20088 17604 20116 17632
rect 17770 17592 17776 17604
rect 10735 17564 11744 17592
rect 13202 17564 17776 17592
rect 10735 17561 10747 17564
rect 10689 17555 10747 17561
rect 4172 17496 6914 17524
rect 7561 17527 7619 17533
rect 3108 17487 3157 17493
rect 7561 17493 7573 17527
rect 7607 17524 7619 17527
rect 7926 17524 7932 17536
rect 7607 17496 7932 17524
rect 7607 17493 7619 17496
rect 7561 17487 7619 17493
rect 3108 17484 3114 17487
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 11716 17524 11744 17564
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 19794 17552 19800 17604
rect 19852 17592 19858 17604
rect 19889 17595 19947 17601
rect 19889 17592 19901 17595
rect 19852 17564 19901 17592
rect 19852 17552 19858 17564
rect 19889 17561 19901 17564
rect 19935 17561 19947 17595
rect 20070 17592 20076 17604
rect 20031 17564 20076 17592
rect 19889 17555 19947 17561
rect 20070 17552 20076 17564
rect 20128 17552 20134 17604
rect 17862 17524 17868 17536
rect 11716 17496 17868 17524
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 17957 17527 18015 17533
rect 17957 17493 17969 17527
rect 18003 17524 18015 17527
rect 18598 17524 18604 17536
rect 18003 17496 18604 17524
rect 18003 17493 18015 17496
rect 17957 17487 18015 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 1104 17434 20859 17456
rect 1104 17382 5848 17434
rect 5900 17382 5912 17434
rect 5964 17382 5976 17434
rect 6028 17382 6040 17434
rect 6092 17382 6104 17434
rect 6156 17382 10747 17434
rect 10799 17382 10811 17434
rect 10863 17382 10875 17434
rect 10927 17382 10939 17434
rect 10991 17382 11003 17434
rect 11055 17382 15646 17434
rect 15698 17382 15710 17434
rect 15762 17382 15774 17434
rect 15826 17382 15838 17434
rect 15890 17382 15902 17434
rect 15954 17382 20545 17434
rect 20597 17382 20609 17434
rect 20661 17382 20673 17434
rect 20725 17382 20737 17434
rect 20789 17382 20801 17434
rect 20853 17382 20859 17434
rect 1104 17360 20859 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 9674 17320 9680 17332
rect 9635 17292 9680 17320
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 12713 17323 12771 17329
rect 12713 17289 12725 17323
rect 12759 17320 12771 17323
rect 15378 17320 15384 17332
rect 12759 17292 15384 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 15378 17280 15384 17292
rect 15436 17320 15442 17332
rect 16482 17320 16488 17332
rect 15436 17292 16488 17320
rect 15436 17280 15442 17292
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 16991 17323 17049 17329
rect 16991 17289 17003 17323
rect 17037 17320 17049 17323
rect 17586 17320 17592 17332
rect 17037 17292 17592 17320
rect 17037 17289 17049 17292
rect 16991 17283 17049 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 2590 17212 2596 17264
rect 2648 17212 2654 17264
rect 3050 17252 3056 17264
rect 3011 17224 3056 17252
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 3142 17212 3148 17264
rect 3200 17252 3206 17264
rect 3200 17224 3372 17252
rect 3200 17212 3206 17224
rect 3344 17193 3372 17224
rect 18598 17212 18604 17264
rect 18656 17212 18662 17264
rect 3878 17193 3884 17196
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 3856 17187 3884 17193
rect 3856 17153 3868 17187
rect 3856 17147 3884 17153
rect 3878 17144 3884 17147
rect 3936 17144 3942 17196
rect 7282 17184 7288 17196
rect 7243 17156 7288 17184
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 7926 17184 7932 17196
rect 7887 17156 7932 17184
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 9490 17184 9496 17196
rect 9451 17156 9496 17184
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 12526 17184 12532 17196
rect 12487 17156 12532 17184
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 14642 17184 14648 17196
rect 14603 17156 14648 17184
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 16888 17187 16946 17193
rect 16888 17184 16900 17187
rect 16163 17156 16900 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16888 17153 16900 17156
rect 16934 17153 16946 17187
rect 17862 17184 17868 17196
rect 17823 17156 17868 17184
rect 16888 17147 16946 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 15470 17116 15476 17128
rect 15335 17088 15476 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 15470 17076 15476 17088
rect 15528 17116 15534 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15528 17088 15945 17116
rect 15528 17076 15534 17088
rect 15933 17085 15945 17088
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17552 17088 18153 17116
rect 17552 17076 17558 17088
rect 18141 17085 18153 17088
rect 18187 17116 18199 17119
rect 18506 17116 18512 17128
rect 18187 17088 18512 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 15749 17051 15807 17057
rect 15749 17017 15761 17051
rect 15795 17048 15807 17051
rect 16022 17048 16028 17060
rect 15795 17020 16028 17048
rect 15795 17017 15807 17020
rect 15749 17011 15807 17017
rect 16022 17008 16028 17020
rect 16080 17008 16086 17060
rect 3970 16989 3976 16992
rect 3927 16983 3976 16989
rect 3927 16949 3939 16983
rect 3973 16949 3976 16983
rect 3927 16943 3976 16949
rect 3970 16940 3976 16943
rect 4028 16940 4034 16992
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 7101 16983 7159 16989
rect 7101 16980 7113 16983
rect 6880 16952 7113 16980
rect 6880 16940 6886 16952
rect 7101 16949 7113 16952
rect 7147 16949 7159 16983
rect 7742 16980 7748 16992
rect 7703 16952 7748 16980
rect 7101 16943 7159 16949
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 19613 16983 19671 16989
rect 19613 16949 19625 16983
rect 19659 16980 19671 16983
rect 19886 16980 19892 16992
rect 19659 16952 19892 16980
rect 19659 16949 19671 16952
rect 19613 16943 19671 16949
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 1104 16890 20700 16912
rect 1104 16838 3399 16890
rect 3451 16838 3463 16890
rect 3515 16838 3527 16890
rect 3579 16838 3591 16890
rect 3643 16838 3655 16890
rect 3707 16838 8298 16890
rect 8350 16838 8362 16890
rect 8414 16838 8426 16890
rect 8478 16838 8490 16890
rect 8542 16838 8554 16890
rect 8606 16838 13197 16890
rect 13249 16838 13261 16890
rect 13313 16838 13325 16890
rect 13377 16838 13389 16890
rect 13441 16838 13453 16890
rect 13505 16838 18096 16890
rect 18148 16838 18160 16890
rect 18212 16838 18224 16890
rect 18276 16838 18288 16890
rect 18340 16838 18352 16890
rect 18404 16838 20700 16890
rect 1104 16816 20700 16838
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 8662 16776 8668 16788
rect 8619 16748 8668 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 8662 16736 8668 16748
rect 8720 16776 8726 16788
rect 9490 16776 9496 16788
rect 8720 16748 9496 16776
rect 8720 16736 8726 16748
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 12526 16776 12532 16788
rect 12483 16748 12532 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 16022 16776 16028 16788
rect 13648 16748 15884 16776
rect 15983 16748 16028 16776
rect 3007 16711 3065 16717
rect 3007 16708 3019 16711
rect 2332 16680 3019 16708
rect 2038 16600 2044 16652
rect 2096 16640 2102 16652
rect 2133 16643 2191 16649
rect 2133 16640 2145 16643
rect 2096 16612 2145 16640
rect 2096 16600 2102 16612
rect 2133 16609 2145 16612
rect 2179 16609 2191 16643
rect 2133 16603 2191 16609
rect 2332 16581 2360 16680
rect 3007 16677 3019 16680
rect 3053 16677 3065 16711
rect 3007 16671 3065 16677
rect 2498 16640 2504 16652
rect 2459 16612 2504 16640
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 3970 16640 3976 16652
rect 3931 16612 3976 16640
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 4522 16640 4528 16652
rect 4172 16612 4528 16640
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 3110 16575 3168 16581
rect 3110 16541 3122 16575
rect 3156 16572 3168 16575
rect 3878 16572 3884 16584
rect 3156 16544 3884 16572
rect 3156 16541 3168 16544
rect 3110 16535 3168 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4172 16581 4200 16612
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7742 16640 7748 16652
rect 7147 16612 7748 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16640 10379 16643
rect 10410 16640 10416 16652
rect 10367 16612 10416 16640
rect 10367 16609 10379 16612
rect 10321 16603 10379 16609
rect 10410 16600 10416 16612
rect 10468 16640 10474 16652
rect 10468 16612 11560 16640
rect 10468 16600 10474 16612
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16574 4215 16575
rect 4341 16575 4399 16581
rect 4203 16546 4237 16574
rect 4203 16541 4215 16546
rect 4157 16535 4215 16541
rect 4341 16541 4353 16575
rect 4387 16572 4399 16575
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 4387 16544 4813 16572
rect 4387 16541 4399 16544
rect 4341 16535 4399 16541
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 10042 16572 10048 16584
rect 10003 16544 10048 16572
rect 4801 16535 4859 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 11532 16572 11560 16612
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 12492 16612 13461 16640
rect 12492 16600 12498 16612
rect 13449 16609 13461 16612
rect 13495 16640 13507 16643
rect 13648 16640 13676 16748
rect 15856 16708 15884 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 15856 16680 16620 16708
rect 13495 16612 13676 16640
rect 13725 16643 13783 16649
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 13771 16612 14565 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 16482 16640 16488 16652
rect 16443 16612 16488 16640
rect 14553 16603 14611 16609
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 16592 16640 16620 16680
rect 16761 16643 16819 16649
rect 16761 16640 16773 16643
rect 16592 16612 16773 16640
rect 16761 16609 16773 16612
rect 16807 16640 16819 16643
rect 17494 16640 17500 16652
rect 16807 16612 17500 16640
rect 16807 16609 16819 16612
rect 16761 16603 16819 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11532 16544 12265 16572
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 13357 16575 13415 16581
rect 13357 16541 13369 16575
rect 13403 16572 13415 16575
rect 14274 16572 14280 16584
rect 13403 16544 13768 16572
rect 14235 16544 14280 16572
rect 13403 16541 13415 16544
rect 13357 16535 13415 16541
rect 13740 16516 13768 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 20162 16572 20168 16584
rect 20123 16544 20168 16572
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 8110 16464 8116 16516
rect 8168 16464 8174 16516
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 9824 16476 10810 16504
rect 9824 16464 9830 16476
rect 13722 16464 13728 16516
rect 13780 16464 13786 16516
rect 15930 16504 15936 16516
rect 15778 16476 15936 16504
rect 15930 16464 15936 16476
rect 15988 16504 15994 16516
rect 16114 16504 16120 16516
rect 15988 16476 16120 16504
rect 15988 16464 15994 16476
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 17770 16464 17776 16516
rect 17828 16464 17834 16516
rect 4985 16439 5043 16445
rect 4985 16405 4997 16439
rect 5031 16436 5043 16439
rect 5626 16436 5632 16448
rect 5031 16408 5632 16436
rect 5031 16405 5043 16408
rect 4985 16399 5043 16405
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 11606 16396 11612 16448
rect 11664 16436 11670 16448
rect 11793 16439 11851 16445
rect 11793 16436 11805 16439
rect 11664 16408 11805 16436
rect 11664 16396 11670 16408
rect 11793 16405 11805 16408
rect 11839 16405 11851 16439
rect 11793 16399 11851 16405
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 18506 16436 18512 16448
rect 18279 16408 18512 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 19978 16436 19984 16448
rect 19939 16408 19984 16436
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 1104 16346 20859 16368
rect 1104 16294 5848 16346
rect 5900 16294 5912 16346
rect 5964 16294 5976 16346
rect 6028 16294 6040 16346
rect 6092 16294 6104 16346
rect 6156 16294 10747 16346
rect 10799 16294 10811 16346
rect 10863 16294 10875 16346
rect 10927 16294 10939 16346
rect 10991 16294 11003 16346
rect 11055 16294 15646 16346
rect 15698 16294 15710 16346
rect 15762 16294 15774 16346
rect 15826 16294 15838 16346
rect 15890 16294 15902 16346
rect 15954 16294 20545 16346
rect 20597 16294 20609 16346
rect 20661 16294 20673 16346
rect 20725 16294 20737 16346
rect 20789 16294 20801 16346
rect 20853 16294 20859 16346
rect 1104 16272 20859 16294
rect 2590 16192 2596 16244
rect 2648 16232 2654 16244
rect 2648 16204 3050 16232
rect 2648 16192 2654 16204
rect 3022 16164 3050 16204
rect 3234 16192 3240 16244
rect 3292 16232 3298 16244
rect 3375 16235 3433 16241
rect 3375 16232 3387 16235
rect 3292 16204 3387 16232
rect 3292 16192 3298 16204
rect 3375 16201 3387 16204
rect 3421 16201 3433 16235
rect 3375 16195 3433 16201
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 7282 16232 7288 16244
rect 7239 16204 7288 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10100 16204 10609 16232
rect 10100 16192 10106 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 14642 16232 14648 16244
rect 14599 16204 14648 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16232 20223 16235
rect 20254 16232 20260 16244
rect 20211 16204 20260 16232
rect 20211 16201 20223 16204
rect 20165 16195 20223 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 3786 16164 3792 16176
rect 2990 16136 3792 16164
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 1627 16068 2084 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1946 16028 1952 16040
rect 1907 16000 1952 16028
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2056 16028 2084 16068
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 6880 16068 7021 16096
rect 6880 16056 6886 16068
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7300 16096 7328 16192
rect 8662 16164 8668 16176
rect 8623 16136 8668 16164
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 17129 16167 17187 16173
rect 17129 16133 17141 16167
rect 17175 16164 17187 16167
rect 17770 16164 17776 16176
rect 17175 16136 17776 16164
rect 17175 16133 17187 16136
rect 17129 16127 17187 16133
rect 17770 16124 17776 16136
rect 17828 16124 17834 16176
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7300 16068 7665 16096
rect 7009 16059 7067 16065
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 9766 16056 9772 16108
rect 9824 16056 9830 16108
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 10560 16068 10793 16096
rect 10560 16056 10566 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11664 16068 12173 16096
rect 11664 16056 11670 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12805 16099 12863 16105
rect 12805 16096 12817 16099
rect 12161 16059 12219 16065
rect 12360 16068 12817 16096
rect 2498 16028 2504 16040
rect 2056 16000 2504 16028
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10410 16028 10416 16040
rect 10183 16000 10416 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 7837 15963 7895 15969
rect 7837 15929 7849 15963
rect 7883 15960 7895 15963
rect 8404 15960 8432 15991
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 12360 15969 12388 16068
rect 12805 16065 12817 16068
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16096 13967 16099
rect 14274 16096 14280 16108
rect 13955 16068 14280 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 7883 15932 8432 15960
rect 12345 15963 12403 15969
rect 7883 15929 7895 15932
rect 7837 15923 7895 15929
rect 12345 15929 12357 15963
rect 12391 15929 12403 15963
rect 12345 15923 12403 15929
rect 12989 15963 13047 15969
rect 12989 15929 13001 15963
rect 13035 15960 13047 15963
rect 13924 15960 13952 16059
rect 14274 16056 14280 16068
rect 14332 16096 14338 16108
rect 15102 16096 15108 16108
rect 14332 16068 15108 16096
rect 14332 16056 14338 16068
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 15470 16096 15476 16108
rect 15431 16068 15476 16096
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 16022 16056 16028 16108
rect 16080 16096 16086 16108
rect 16234 16099 16292 16105
rect 16234 16096 16246 16099
rect 16080 16068 16246 16096
rect 16080 16056 16086 16068
rect 16234 16065 16246 16068
rect 16280 16065 16292 16099
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 16234 16059 16292 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 17736 16068 17954 16096
rect 17736 16056 17742 16068
rect 17926 16028 17954 16068
rect 19794 16056 19800 16108
rect 19852 16056 19858 16108
rect 18414 16028 18420 16040
rect 17926 16000 18420 16028
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 13035 15932 13952 15960
rect 15657 15963 15715 15969
rect 13035 15929 13047 15932
rect 12989 15923 13047 15929
rect 15657 15929 15669 15963
rect 15703 15960 15715 15963
rect 16163 15963 16221 15969
rect 16163 15960 16175 15963
rect 15703 15932 16175 15960
rect 15703 15929 15715 15932
rect 15657 15923 15715 15929
rect 16163 15929 16175 15932
rect 16209 15929 16221 15963
rect 16163 15923 16221 15929
rect 1104 15802 20700 15824
rect 1104 15750 3399 15802
rect 3451 15750 3463 15802
rect 3515 15750 3527 15802
rect 3579 15750 3591 15802
rect 3643 15750 3655 15802
rect 3707 15750 8298 15802
rect 8350 15750 8362 15802
rect 8414 15750 8426 15802
rect 8478 15750 8490 15802
rect 8542 15750 8554 15802
rect 8606 15750 13197 15802
rect 13249 15750 13261 15802
rect 13313 15750 13325 15802
rect 13377 15750 13389 15802
rect 13441 15750 13453 15802
rect 13505 15750 18096 15802
rect 18148 15750 18160 15802
rect 18212 15750 18224 15802
rect 18276 15750 18288 15802
rect 18340 15750 18352 15802
rect 18404 15750 20700 15802
rect 1104 15728 20700 15750
rect 1946 15697 1952 15700
rect 1903 15691 1952 15697
rect 1903 15657 1915 15691
rect 1949 15657 1952 15691
rect 1903 15651 1952 15657
rect 1946 15648 1952 15651
rect 2004 15648 2010 15700
rect 17313 15691 17371 15697
rect 17313 15657 17325 15691
rect 17359 15688 17371 15691
rect 18690 15688 18696 15700
rect 17359 15660 18696 15688
rect 17359 15657 17371 15660
rect 17313 15651 17371 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 7653 15623 7711 15629
rect 7653 15589 7665 15623
rect 7699 15589 7711 15623
rect 7653 15583 7711 15589
rect 10045 15623 10103 15629
rect 10045 15589 10057 15623
rect 10091 15620 10103 15623
rect 10091 15592 10640 15620
rect 10091 15589 10103 15592
rect 10045 15583 10103 15589
rect 1486 15444 1492 15496
rect 1544 15484 1550 15496
rect 2006 15487 2064 15493
rect 2006 15484 2018 15487
rect 1544 15456 2018 15484
rect 1544 15444 1550 15456
rect 2006 15453 2018 15456
rect 2052 15484 2064 15487
rect 2682 15484 2688 15496
rect 2052 15456 2688 15484
rect 2052 15453 2064 15456
rect 2006 15447 2064 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 6880 15456 7481 15484
rect 6880 15444 6886 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7668 15484 7696 15583
rect 10612 15561 10640 15592
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 13780 15592 15240 15620
rect 13780 15580 13786 15592
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 11606 15552 11612 15564
rect 10919 15524 11612 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 15102 15552 15108 15564
rect 15063 15524 15108 15552
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 15212 15552 15240 15592
rect 17034 15580 17040 15632
rect 17092 15620 17098 15632
rect 18325 15623 18383 15629
rect 18325 15620 18337 15623
rect 17092 15592 18337 15620
rect 17092 15580 17098 15592
rect 18325 15589 18337 15592
rect 18371 15589 18383 15623
rect 18325 15583 18383 15589
rect 17586 15552 17592 15564
rect 15212 15524 17592 15552
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 7668 15456 9873 15484
rect 7469 15447 7527 15453
rect 9861 15453 9873 15456
rect 9907 15484 9919 15487
rect 10502 15484 10508 15496
rect 9907 15456 10508 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 18506 15444 18512 15496
rect 18564 15444 18570 15496
rect 20070 15484 20076 15496
rect 20031 15456 20076 15484
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 7282 15376 7288 15428
rect 7340 15416 7346 15428
rect 8110 15416 8116 15428
rect 7340 15388 8116 15416
rect 7340 15376 7346 15388
rect 8110 15376 8116 15388
rect 8168 15416 8174 15428
rect 9766 15416 9772 15428
rect 8168 15388 9772 15416
rect 8168 15376 8174 15388
rect 9766 15376 9772 15388
rect 9824 15416 9830 15428
rect 9824 15388 11362 15416
rect 9824 15376 9830 15388
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 15381 15419 15439 15425
rect 15381 15416 15393 15419
rect 14148 15388 15393 15416
rect 14148 15376 14154 15388
rect 15381 15385 15393 15388
rect 15427 15385 15439 15419
rect 15381 15379 15439 15385
rect 16114 15376 16120 15428
rect 16172 15376 16178 15428
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 19392 15388 19717 15416
rect 19392 15376 19398 15388
rect 19705 15385 19717 15388
rect 19751 15385 19763 15419
rect 19705 15379 19763 15385
rect 12342 15348 12348 15360
rect 12303 15320 12348 15348
rect 12342 15308 12348 15320
rect 12400 15308 12406 15360
rect 16850 15348 16856 15360
rect 16811 15320 16856 15348
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 18690 15348 18696 15360
rect 18651 15320 18696 15348
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 1104 15258 20859 15280
rect 1104 15206 5848 15258
rect 5900 15206 5912 15258
rect 5964 15206 5976 15258
rect 6028 15206 6040 15258
rect 6092 15206 6104 15258
rect 6156 15206 10747 15258
rect 10799 15206 10811 15258
rect 10863 15206 10875 15258
rect 10927 15206 10939 15258
rect 10991 15206 11003 15258
rect 11055 15206 15646 15258
rect 15698 15206 15710 15258
rect 15762 15206 15774 15258
rect 15826 15206 15838 15258
rect 15890 15206 15902 15258
rect 15954 15206 20545 15258
rect 20597 15206 20609 15258
rect 20661 15206 20673 15258
rect 20725 15206 20737 15258
rect 20789 15206 20801 15258
rect 20853 15206 20859 15258
rect 1104 15184 20859 15206
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 9582 15144 9588 15156
rect 8168 15116 9588 15144
rect 8168 15104 8174 15116
rect 9582 15104 9588 15116
rect 9640 15144 9646 15156
rect 12894 15144 12900 15156
rect 9640 15116 12900 15144
rect 9640 15104 9646 15116
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 20162 15144 20168 15156
rect 20123 15116 20168 15144
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 5626 15036 5632 15088
rect 5684 15076 5690 15088
rect 18690 15076 18696 15088
rect 5684 15048 7512 15076
rect 18651 15048 18696 15076
rect 5684 15036 5690 15048
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 5350 15008 5356 15020
rect 5311 14980 5356 15008
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 7484 15017 7512 15048
rect 18690 15036 18696 15048
rect 18748 15036 18754 15088
rect 19334 15036 19340 15088
rect 19392 15036 19398 15088
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 10388 15011 10446 15017
rect 10388 14977 10400 15011
rect 10434 15008 10446 15011
rect 10870 15008 10876 15020
rect 10434 14980 10876 15008
rect 10434 14977 10446 14980
rect 10388 14971 10446 14977
rect 6932 14872 6960 14971
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9232 14940 9260 14971
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11977 15011 12035 15017
rect 11977 15008 11989 15011
rect 11204 14980 11989 15008
rect 11204 14968 11210 14980
rect 11977 14977 11989 14980
rect 12023 15008 12035 15011
rect 12342 15008 12348 15020
rect 12023 14980 12348 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 14090 15017 14096 15020
rect 14068 15011 14096 15017
rect 14068 14977 14080 15011
rect 14068 14971 14096 14977
rect 14090 14968 14096 14971
rect 14148 14968 14154 15020
rect 16482 14940 16488 14952
rect 9180 14912 16488 14940
rect 9180 14900 9186 14912
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 18414 14940 18420 14952
rect 18327 14912 18420 14940
rect 18414 14900 18420 14912
rect 18472 14940 18478 14952
rect 18782 14940 18788 14952
rect 18472 14912 18788 14940
rect 18472 14900 18478 14912
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 7558 14872 7564 14884
rect 6932 14844 7564 14872
rect 7558 14832 7564 14844
rect 7616 14872 7622 14884
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 7616 14844 7665 14872
rect 7616 14832 7622 14844
rect 7653 14841 7665 14844
rect 7699 14841 7711 14875
rect 7653 14835 7711 14841
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14804 1823 14807
rect 1854 14804 1860 14816
rect 1811 14776 1860 14804
rect 1811 14773 1823 14776
rect 1765 14767 1823 14773
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14804 6883 14807
rect 7282 14804 7288 14816
rect 6871 14776 7288 14804
rect 6871 14773 6883 14776
rect 6825 14767 6883 14773
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 9950 14804 9956 14816
rect 9907 14776 9956 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10459 14807 10517 14813
rect 10459 14773 10471 14807
rect 10505 14804 10517 14807
rect 11330 14804 11336 14816
rect 10505 14776 11336 14804
rect 10505 14773 10517 14776
rect 10459 14767 10517 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 12161 14807 12219 14813
rect 12161 14773 12173 14807
rect 12207 14804 12219 14807
rect 12250 14804 12256 14816
rect 12207 14776 12256 14804
rect 12207 14773 12219 14776
rect 12161 14767 12219 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 14139 14807 14197 14813
rect 14139 14773 14151 14807
rect 14185 14804 14197 14807
rect 14550 14804 14556 14816
rect 14185 14776 14556 14804
rect 14185 14773 14197 14776
rect 14139 14767 14197 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 1104 14714 20700 14736
rect 1104 14662 3399 14714
rect 3451 14662 3463 14714
rect 3515 14662 3527 14714
rect 3579 14662 3591 14714
rect 3643 14662 3655 14714
rect 3707 14662 8298 14714
rect 8350 14662 8362 14714
rect 8414 14662 8426 14714
rect 8478 14662 8490 14714
rect 8542 14662 8554 14714
rect 8606 14662 13197 14714
rect 13249 14662 13261 14714
rect 13313 14662 13325 14714
rect 13377 14662 13389 14714
rect 13441 14662 13453 14714
rect 13505 14662 18096 14714
rect 18148 14662 18160 14714
rect 18212 14662 18224 14714
rect 18276 14662 18288 14714
rect 18340 14662 18352 14714
rect 18404 14662 20700 14714
rect 1104 14640 20700 14662
rect 6886 14572 10548 14600
rect 4893 14535 4951 14541
rect 4893 14501 4905 14535
rect 4939 14532 4951 14535
rect 4939 14504 5396 14532
rect 4939 14501 4951 14504
rect 4893 14495 4951 14501
rect 5368 14473 5396 14504
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 6886 14464 6914 14572
rect 7929 14535 7987 14541
rect 7929 14501 7941 14535
rect 7975 14501 7987 14535
rect 10520 14532 10548 14572
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 10870 14600 10876 14612
rect 10652 14572 10876 14600
rect 10652 14560 10658 14572
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 13081 14603 13139 14609
rect 13081 14569 13093 14603
rect 13127 14600 13139 14603
rect 14090 14600 14096 14612
rect 13127 14572 14096 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 16025 14603 16083 14609
rect 16025 14569 16037 14603
rect 16071 14600 16083 14603
rect 16574 14600 16580 14612
rect 16071 14572 16580 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17034 14600 17040 14612
rect 16995 14572 17040 14600
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 11146 14532 11152 14544
rect 10520 14504 11152 14532
rect 7929 14495 7987 14501
rect 5675 14436 6914 14464
rect 7944 14464 7972 14495
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 11330 14532 11336 14544
rect 11291 14504 11336 14532
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 17402 14492 17408 14544
rect 17460 14532 17466 14544
rect 18049 14535 18107 14541
rect 18049 14532 18061 14535
rect 17460 14504 18061 14532
rect 17460 14492 17466 14504
rect 18049 14501 18061 14504
rect 18095 14501 18107 14535
rect 18049 14495 18107 14501
rect 9122 14464 9128 14476
rect 7944 14436 9128 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 9122 14424 9128 14436
rect 9180 14424 9186 14476
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 10468 14436 11529 14464
rect 10468 14424 10474 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 14550 14464 14556 14476
rect 14511 14436 14556 14464
rect 11517 14427 11575 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 17586 14424 17592 14476
rect 17644 14424 17650 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1854 14396 1860 14408
rect 1719 14368 1860 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 4755 14368 5396 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 5368 14340 5396 14368
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7432 14368 7757 14396
rect 7432 14356 7438 14368
rect 7745 14365 7757 14368
rect 7791 14365 7803 14399
rect 12250 14396 12256 14408
rect 12211 14368 12256 14396
rect 7745 14359 7803 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 12894 14396 12900 14408
rect 12855 14368 12900 14396
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 16908 14368 17250 14396
rect 16908 14356 16914 14368
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 4522 14328 4528 14340
rect 2823 14300 4528 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 4522 14288 4528 14300
rect 4580 14288 4586 14340
rect 5350 14288 5356 14340
rect 5408 14288 5414 14340
rect 7282 14328 7288 14340
rect 6854 14300 7288 14328
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 8754 14288 8760 14340
rect 8812 14328 8818 14340
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 8812 14300 9413 14328
rect 8812 14288 8818 14300
rect 9401 14297 9413 14300
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 9858 14288 9864 14340
rect 9916 14288 9922 14340
rect 12437 14331 12495 14337
rect 12437 14297 12449 14331
rect 12483 14328 12495 14331
rect 12526 14328 12532 14340
rect 12483 14300 12532 14328
rect 12483 14297 12495 14300
rect 12437 14291 12495 14297
rect 12526 14288 12532 14300
rect 12584 14328 12590 14340
rect 14292 14328 14320 14356
rect 12584 14300 14320 14328
rect 12584 14288 12590 14300
rect 15194 14288 15200 14340
rect 15252 14288 15258 14340
rect 1857 14263 1915 14269
rect 1857 14229 1869 14263
rect 1903 14260 1915 14263
rect 1946 14260 1952 14272
rect 1903 14232 1952 14260
rect 1903 14229 1915 14232
rect 1857 14223 1915 14229
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 2685 14263 2743 14269
rect 2685 14229 2697 14263
rect 2731 14260 2743 14263
rect 2866 14260 2872 14272
rect 2731 14232 2872 14260
rect 2731 14229 2743 14232
rect 2685 14223 2743 14229
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 7101 14263 7159 14269
rect 7101 14229 7113 14263
rect 7147 14260 7159 14263
rect 7190 14260 7196 14272
rect 7147 14232 7196 14260
rect 7147 14229 7159 14232
rect 7101 14223 7159 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 11514 14220 11520 14272
rect 11572 14260 11578 14272
rect 11698 14260 11704 14272
rect 11572 14232 11704 14260
rect 11572 14220 11578 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 18414 14260 18420 14272
rect 18375 14232 18420 14260
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 1104 14170 20859 14192
rect 1104 14118 5848 14170
rect 5900 14118 5912 14170
rect 5964 14118 5976 14170
rect 6028 14118 6040 14170
rect 6092 14118 6104 14170
rect 6156 14118 10747 14170
rect 10799 14118 10811 14170
rect 10863 14118 10875 14170
rect 10927 14118 10939 14170
rect 10991 14118 11003 14170
rect 11055 14118 15646 14170
rect 15698 14118 15710 14170
rect 15762 14118 15774 14170
rect 15826 14118 15838 14170
rect 15890 14118 15902 14170
rect 15954 14118 20545 14170
rect 20597 14118 20609 14170
rect 20661 14118 20673 14170
rect 20725 14118 20737 14170
rect 20789 14118 20801 14170
rect 20853 14118 20859 14170
rect 1104 14096 20859 14118
rect 4062 14065 4068 14068
rect 4019 14059 4068 14065
rect 4019 14025 4031 14059
rect 4065 14025 4068 14059
rect 4019 14019 4068 14025
rect 4062 14016 4068 14019
rect 4120 14016 4126 14068
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 5537 14059 5595 14065
rect 5537 14056 5549 14059
rect 5408 14028 5549 14056
rect 5408 14016 5414 14028
rect 5537 14025 5549 14028
rect 5583 14025 5595 14059
rect 7374 14056 7380 14068
rect 7335 14028 7380 14056
rect 5537 14019 5595 14025
rect 7374 14016 7380 14028
rect 7432 14016 7438 14068
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10468 14028 10609 14056
rect 10468 14016 10474 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 10597 14019 10655 14025
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14056 14335 14059
rect 14366 14056 14372 14068
rect 14323 14028 14372 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 3786 13988 3792 14000
rect 3634 13960 3792 13988
rect 3786 13948 3792 13960
rect 3844 13988 3850 14000
rect 9858 13988 9864 14000
rect 3844 13960 9864 13988
rect 3844 13948 3850 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 14642 13988 14648 14000
rect 14030 13960 14648 13988
rect 14642 13948 14648 13960
rect 14700 13948 14706 14000
rect 18414 13948 18420 14000
rect 18472 13988 18478 14000
rect 18693 13991 18751 13997
rect 18693 13988 18705 13991
rect 18472 13960 18705 13988
rect 18472 13948 18478 13960
rect 18693 13957 18705 13960
rect 18739 13957 18751 13991
rect 18693 13951 18751 13957
rect 19334 13948 19340 14000
rect 19392 13948 19398 14000
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1616 13923 1674 13929
rect 1616 13920 1628 13923
rect 1544 13892 1628 13920
rect 1544 13880 1550 13892
rect 1616 13889 1628 13892
rect 1662 13889 1674 13923
rect 1616 13883 1674 13889
rect 1719 13923 1777 13929
rect 1719 13889 1731 13923
rect 1765 13920 1777 13923
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 1765 13892 2605 13920
rect 1765 13889 1777 13892
rect 1719 13883 1777 13889
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 4706 13920 4712 13932
rect 4667 13892 4712 13920
rect 2593 13883 2651 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 6822 13920 6828 13932
rect 5767 13892 6828 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 7190 13920 7196 13932
rect 7151 13892 7196 13920
rect 7190 13880 7196 13892
rect 7248 13880 7254 13932
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8260 13892 8401 13920
rect 8260 13880 8266 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 9950 13920 9956 13932
rect 9911 13892 9956 13920
rect 8389 13883 8447 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11736 13923 11794 13929
rect 11736 13920 11748 13923
rect 11112 13892 11748 13920
rect 11112 13880 11118 13892
rect 11736 13889 11748 13892
rect 11782 13889 11794 13923
rect 12526 13920 12532 13932
rect 12487 13892 12532 13920
rect 11736 13883 11794 13889
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 6454 13852 6460 13864
rect 2271 13824 6460 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 8168 13824 8309 13852
rect 8168 13812 8174 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8297 13815 8355 13821
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 11839 13855 11897 13861
rect 11839 13821 11851 13855
rect 11885 13852 11897 13855
rect 12434 13852 12440 13864
rect 11885 13824 12440 13852
rect 11885 13821 11897 13824
rect 11839 13815 11897 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13852 18475 13855
rect 18782 13852 18788 13864
rect 18463 13824 18788 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 20162 13716 20168 13728
rect 20123 13688 20168 13716
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 1104 13626 20700 13648
rect 1104 13574 3399 13626
rect 3451 13574 3463 13626
rect 3515 13574 3527 13626
rect 3579 13574 3591 13626
rect 3643 13574 3655 13626
rect 3707 13574 8298 13626
rect 8350 13574 8362 13626
rect 8414 13574 8426 13626
rect 8478 13574 8490 13626
rect 8542 13574 8554 13626
rect 8606 13574 13197 13626
rect 13249 13574 13261 13626
rect 13313 13574 13325 13626
rect 13377 13574 13389 13626
rect 13441 13574 13453 13626
rect 13505 13574 18096 13626
rect 18148 13574 18160 13626
rect 18212 13574 18224 13626
rect 18276 13574 18288 13626
rect 18340 13574 18352 13626
rect 18404 13574 20700 13626
rect 1104 13552 20700 13574
rect 2133 13515 2191 13521
rect 2133 13481 2145 13515
rect 2179 13512 2191 13515
rect 4706 13512 4712 13524
rect 2179 13484 4712 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 11054 13512 11060 13524
rect 11015 13484 11060 13512
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13311 13515 13369 13521
rect 13311 13512 13323 13515
rect 12860 13484 13323 13512
rect 12860 13472 12866 13484
rect 13311 13481 13323 13484
rect 13357 13481 13369 13515
rect 13311 13475 13369 13481
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 14090 13512 14096 13524
rect 13504 13484 14096 13512
rect 13504 13472 13510 13484
rect 14090 13472 14096 13484
rect 14148 13512 14154 13524
rect 14534 13515 14592 13521
rect 14534 13512 14546 13515
rect 14148 13484 14546 13512
rect 14148 13472 14154 13484
rect 14534 13481 14546 13484
rect 14580 13512 14592 13515
rect 19978 13512 19984 13524
rect 14580 13484 15976 13512
rect 19939 13484 19984 13512
rect 14580 13481 14592 13484
rect 14534 13475 14592 13481
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 2685 13447 2743 13453
rect 2685 13444 2697 13447
rect 1544 13416 2697 13444
rect 1544 13404 1550 13416
rect 2685 13413 2697 13416
rect 2731 13413 2743 13447
rect 2685 13407 2743 13413
rect 10594 13404 10600 13456
rect 10652 13444 10658 13456
rect 10689 13447 10747 13453
rect 10689 13444 10701 13447
rect 10652 13416 10701 13444
rect 10652 13404 10658 13416
rect 10689 13413 10701 13416
rect 10735 13413 10747 13447
rect 10689 13407 10747 13413
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 12492 13416 12537 13444
rect 12492 13404 12498 13416
rect 5534 13376 5540 13388
rect 5495 13348 5540 13376
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 7190 13376 7196 13388
rect 5859 13348 7196 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 10468 13348 10885 13376
rect 10468 13336 10474 13348
rect 10873 13345 10885 13348
rect 10919 13345 10931 13379
rect 10873 13339 10931 13345
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 15194 13376 15200 13388
rect 12851 13348 15200 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15948 13376 15976 13484
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 15948 13348 16773 13376
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 1946 13308 1952 13320
rect 1907 13280 1952 13308
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 2866 13308 2872 13320
rect 2779 13280 2872 13308
rect 2866 13268 2872 13280
rect 2924 13308 2930 13320
rect 4522 13308 4528 13320
rect 2924 13280 4528 13308
rect 2924 13268 2930 13280
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 12618 13308 12624 13320
rect 12579 13280 12624 13308
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13446 13317 13452 13320
rect 13414 13311 13452 13317
rect 13414 13308 13426 13311
rect 13136 13280 13426 13308
rect 13136 13268 13142 13280
rect 13414 13277 13426 13280
rect 13414 13271 13452 13277
rect 13446 13268 13452 13271
rect 13504 13268 13510 13320
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14274 13308 14280 13320
rect 13964 13280 14280 13308
rect 13964 13268 13970 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 16482 13308 16488 13320
rect 16443 13280 16488 13308
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 20162 13308 20168 13320
rect 20123 13280 20168 13308
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 7300 13240 7328 13268
rect 7742 13240 7748 13252
rect 7038 13212 7748 13240
rect 7742 13200 7748 13212
rect 7800 13200 7806 13252
rect 15194 13200 15200 13252
rect 15252 13200 15258 13252
rect 16114 13200 16120 13252
rect 16172 13240 16178 13252
rect 16172 13212 17250 13240
rect 16172 13200 16178 13212
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 7156 13144 7297 13172
rect 7156 13132 7162 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 7285 13135 7343 13141
rect 16025 13175 16083 13181
rect 16025 13141 16037 13175
rect 16071 13172 16083 13175
rect 16666 13172 16672 13184
rect 16071 13144 16672 13172
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18598 13172 18604 13184
rect 18279 13144 18604 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 1104 13082 20859 13104
rect 1104 13030 5848 13082
rect 5900 13030 5912 13082
rect 5964 13030 5976 13082
rect 6028 13030 6040 13082
rect 6092 13030 6104 13082
rect 6156 13030 10747 13082
rect 10799 13030 10811 13082
rect 10863 13030 10875 13082
rect 10927 13030 10939 13082
rect 10991 13030 11003 13082
rect 11055 13030 15646 13082
rect 15698 13030 15710 13082
rect 15762 13030 15774 13082
rect 15826 13030 15838 13082
rect 15890 13030 15902 13082
rect 15954 13030 20545 13082
rect 20597 13030 20609 13082
rect 20661 13030 20673 13082
rect 20725 13030 20737 13082
rect 20789 13030 20801 13082
rect 20853 13030 20859 13082
rect 1104 13008 20859 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12937 2191 12971
rect 2133 12931 2191 12937
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12968 12771 12971
rect 14642 12968 14648 12980
rect 12759 12940 14648 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2038 12832 2044 12844
rect 1995 12804 2044 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2148 12832 2176 12931
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 16117 12971 16175 12977
rect 16117 12968 16129 12971
rect 15028 12940 16129 12968
rect 6825 12903 6883 12909
rect 6825 12869 6837 12903
rect 6871 12900 6883 12903
rect 7098 12900 7104 12912
rect 6871 12872 7104 12900
rect 6871 12869 6883 12872
rect 6825 12863 6883 12869
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 7558 12860 7564 12912
rect 7616 12860 7622 12912
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 15028 12909 15056 12940
rect 16117 12937 16129 12940
rect 16163 12968 16175 12971
rect 16942 12968 16948 12980
rect 16163 12940 16948 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 15013 12903 15071 12909
rect 15013 12900 15025 12903
rect 14148 12872 15025 12900
rect 14148 12860 14154 12872
rect 15013 12869 15025 12872
rect 15059 12869 15071 12903
rect 15013 12863 15071 12869
rect 19334 12860 19340 12912
rect 19392 12860 19398 12912
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2148 12804 2789 12832
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 4338 12832 4344 12844
rect 4299 12804 4344 12832
rect 2777 12795 2835 12801
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 8754 12832 8760 12844
rect 8715 12804 8760 12832
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9950 12832 9956 12844
rect 9911 12804 9956 12832
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 13658 12835 13716 12841
rect 13658 12832 13670 12835
rect 12115 12804 13670 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 13658 12801 13670 12804
rect 13704 12801 13716 12835
rect 13658 12795 13716 12801
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 15620 12804 16221 12832
rect 15620 12792 15626 12804
rect 16209 12801 16221 12804
rect 16255 12832 16267 12835
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 16255 12804 17417 12832
rect 16255 12801 16267 12804
rect 16209 12795 16267 12801
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 6546 12764 6552 12776
rect 6507 12736 6552 12764
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11296 12736 11897 12764
rect 11296 12724 11302 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12676 12736 12909 12764
rect 12676 12724 12682 12736
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 12943 12736 15301 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 15289 12733 15301 12736
rect 15335 12764 15347 12767
rect 16114 12764 16120 12776
rect 15335 12736 16120 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 17681 12767 17739 12773
rect 17681 12733 17693 12767
rect 17727 12764 17739 12767
rect 17770 12764 17776 12776
rect 17727 12736 17776 12764
rect 17727 12733 17739 12736
rect 17681 12727 17739 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 18414 12764 18420 12776
rect 18375 12736 18420 12764
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18690 12764 18696 12776
rect 18651 12736 18696 12764
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 11698 12696 11704 12708
rect 11659 12668 11704 12696
rect 11698 12656 11704 12668
rect 11756 12656 11762 12708
rect 13081 12699 13139 12705
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 13587 12699 13645 12705
rect 13587 12696 13599 12699
rect 13127 12668 13599 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 13587 12665 13599 12668
rect 13633 12665 13645 12699
rect 13587 12659 13645 12665
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 2593 12631 2651 12637
rect 2593 12628 2605 12631
rect 1636 12600 2605 12628
rect 1636 12588 1642 12600
rect 2593 12597 2605 12600
rect 2639 12597 2651 12631
rect 2593 12591 2651 12597
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12628 4583 12631
rect 5166 12628 5172 12640
rect 4571 12600 5172 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 8297 12631 8355 12637
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 8662 12628 8668 12640
rect 8343 12600 8668 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 8941 12631 8999 12637
rect 8941 12597 8953 12631
rect 8987 12628 8999 12631
rect 9122 12628 9128 12640
rect 8987 12600 9128 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 9122 12588 9128 12600
rect 9180 12628 9186 12640
rect 9950 12628 9956 12640
rect 9180 12600 9956 12628
rect 9180 12588 9186 12600
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10502 12588 10508 12640
rect 10560 12628 10566 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10560 12600 10609 12628
rect 10560 12588 10566 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 20162 12628 20168 12640
rect 20123 12600 20168 12628
rect 10597 12591 10655 12597
rect 20162 12588 20168 12600
rect 20220 12588 20226 12640
rect 1104 12538 20700 12560
rect 1104 12486 3399 12538
rect 3451 12486 3463 12538
rect 3515 12486 3527 12538
rect 3579 12486 3591 12538
rect 3643 12486 3655 12538
rect 3707 12486 8298 12538
rect 8350 12486 8362 12538
rect 8414 12486 8426 12538
rect 8478 12486 8490 12538
rect 8542 12486 8554 12538
rect 8606 12486 13197 12538
rect 13249 12486 13261 12538
rect 13313 12486 13325 12538
rect 13377 12486 13389 12538
rect 13441 12486 13453 12538
rect 13505 12486 18096 12538
rect 18148 12486 18160 12538
rect 18212 12486 18224 12538
rect 18276 12486 18288 12538
rect 18340 12486 18352 12538
rect 18404 12486 20700 12538
rect 1104 12464 20700 12486
rect 5997 12427 6055 12433
rect 5997 12393 6009 12427
rect 6043 12424 6055 12427
rect 6546 12424 6552 12436
rect 6043 12396 6552 12424
rect 6043 12393 6055 12396
rect 5997 12387 6055 12393
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 7561 12427 7619 12433
rect 7561 12393 7573 12427
rect 7607 12424 7619 12427
rect 8754 12424 8760 12436
rect 7607 12396 8760 12424
rect 7607 12393 7619 12396
rect 7561 12387 7619 12393
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 10873 12427 10931 12433
rect 10873 12393 10885 12427
rect 10919 12424 10931 12427
rect 11146 12424 11152 12436
rect 10919 12396 11152 12424
rect 10919 12393 10931 12396
rect 10873 12387 10931 12393
rect 11146 12384 11152 12396
rect 11204 12424 11210 12436
rect 11698 12424 11704 12436
rect 11204 12396 11704 12424
rect 11204 12384 11210 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 14182 12424 14188 12436
rect 13495 12396 14188 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 18690 12384 18696 12436
rect 18748 12424 18754 12436
rect 18785 12427 18843 12433
rect 18785 12424 18797 12427
rect 18748 12396 18797 12424
rect 18748 12384 18754 12396
rect 18785 12393 18797 12396
rect 18831 12393 18843 12427
rect 18785 12387 18843 12393
rect 8573 12359 8631 12365
rect 8573 12325 8585 12359
rect 8619 12356 8631 12359
rect 8619 12328 9260 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 8110 12288 8116 12300
rect 8071 12260 8116 12288
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 9122 12288 9128 12300
rect 9083 12260 9128 12288
rect 9122 12248 9128 12260
rect 9180 12248 9186 12300
rect 9232 12288 9260 12328
rect 13078 12316 13084 12368
rect 13136 12356 13142 12368
rect 13136 12328 15332 12356
rect 13136 12316 13142 12328
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 9232 12260 9413 12288
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 15197 12291 15255 12297
rect 15197 12288 15209 12291
rect 10008 12260 15209 12288
rect 10008 12248 10014 12260
rect 15197 12257 15209 12260
rect 15243 12257 15255 12291
rect 15304 12288 15332 12328
rect 18138 12316 18144 12368
rect 18196 12356 18202 12368
rect 18417 12359 18475 12365
rect 18417 12356 18429 12359
rect 18196 12328 18429 12356
rect 18196 12316 18202 12328
rect 18417 12325 18429 12328
rect 18463 12325 18475 12359
rect 19978 12356 19984 12368
rect 19939 12328 19984 12356
rect 18417 12319 18475 12325
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15304 12260 15485 12288
rect 15197 12251 15255 12257
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 18046 12248 18052 12300
rect 18104 12248 18110 12300
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4798 12220 4804 12232
rect 4755 12192 4804 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5166 12220 5172 12232
rect 5127 12192 5172 12220
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12220 5871 12223
rect 6178 12220 6184 12232
rect 5859 12192 6184 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 6178 12180 6184 12192
rect 6236 12220 6242 12232
rect 6641 12223 6699 12229
rect 6236 12192 6500 12220
rect 6236 12180 6242 12192
rect 1762 12084 1768 12096
rect 1723 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 4525 12087 4583 12093
rect 4525 12084 4537 12087
rect 3568 12056 4537 12084
rect 3568 12044 3574 12056
rect 4525 12053 4537 12056
rect 4571 12053 4583 12087
rect 4525 12047 4583 12053
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 6472 12093 6500 12192
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6822 12220 6828 12232
rect 6687 12192 6828 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7156 12192 7389 12220
rect 7156 12180 7162 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 8202 12220 8208 12232
rect 8163 12192 8208 12220
rect 7377 12183 7435 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 14550 12220 14556 12232
rect 14511 12192 14556 12220
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 18598 12180 18604 12232
rect 18656 12180 18662 12232
rect 20162 12220 20168 12232
rect 20123 12192 20168 12220
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 9858 12152 9864 12164
rect 9784 12124 9864 12152
rect 5353 12087 5411 12093
rect 5353 12084 5365 12087
rect 5316 12056 5365 12084
rect 5316 12044 5322 12056
rect 5353 12053 5365 12056
rect 5399 12053 5411 12087
rect 5353 12047 5411 12053
rect 6457 12087 6515 12093
rect 6457 12053 6469 12087
rect 6503 12053 6515 12087
rect 9784 12084 9812 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 11974 12152 11980 12164
rect 11935 12124 11980 12152
rect 11974 12112 11980 12124
rect 12032 12112 12038 12164
rect 12618 12112 12624 12164
rect 12676 12112 12682 12164
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14056 12124 14412 12152
rect 14056 12112 14062 12124
rect 14090 12084 14096 12096
rect 9784 12056 14096 12084
rect 6457 12047 6515 12053
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14384 12093 14412 12124
rect 16114 12112 16120 12164
rect 16172 12112 16178 12164
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12053 14427 12087
rect 16942 12084 16948 12096
rect 16903 12056 16948 12084
rect 14369 12047 14427 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 1104 11994 20859 12016
rect 1104 11942 5848 11994
rect 5900 11942 5912 11994
rect 5964 11942 5976 11994
rect 6028 11942 6040 11994
rect 6092 11942 6104 11994
rect 6156 11942 10747 11994
rect 10799 11942 10811 11994
rect 10863 11942 10875 11994
rect 10927 11942 10939 11994
rect 10991 11942 11003 11994
rect 11055 11942 15646 11994
rect 15698 11942 15710 11994
rect 15762 11942 15774 11994
rect 15826 11942 15838 11994
rect 15890 11942 15902 11994
rect 15954 11942 20545 11994
rect 20597 11942 20609 11994
rect 20661 11942 20673 11994
rect 20725 11942 20737 11994
rect 20789 11942 20801 11994
rect 20853 11942 20859 11994
rect 1104 11920 20859 11942
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 4338 11880 4344 11892
rect 3743 11852 4344 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4798 11880 4804 11892
rect 4759 11852 4804 11880
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 6822 11880 6828 11892
rect 6687 11852 6828 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 11149 11883 11207 11889
rect 11149 11849 11161 11883
rect 11195 11880 11207 11883
rect 11238 11880 11244 11892
rect 11195 11852 11244 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11974 11889 11980 11892
rect 11931 11883 11980 11889
rect 11931 11849 11943 11883
rect 11977 11849 11980 11883
rect 11931 11843 11980 11849
rect 11974 11840 11980 11843
rect 12032 11840 12038 11892
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 18138 11880 18144 11892
rect 16991 11852 18144 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 13906 11812 13912 11824
rect 13648 11784 13912 11812
rect 3510 11744 3516 11756
rect 3471 11716 3516 11744
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4614 11744 4620 11756
rect 4203 11716 4620 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6178 11744 6184 11756
rect 5859 11716 6184 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 6822 11744 6828 11756
rect 6779 11716 6828 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 9928 11747 9986 11753
rect 9928 11713 9940 11747
rect 9974 11744 9986 11747
rect 10502 11744 10508 11756
rect 9974 11716 10364 11744
rect 10463 11716 10508 11744
rect 9974 11713 9986 11716
rect 9928 11707 9986 11713
rect 10336 11676 10364 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 11860 11747 11918 11753
rect 11860 11713 11872 11747
rect 11906 11744 11918 11747
rect 13078 11744 13084 11756
rect 11906 11716 13084 11744
rect 11906 11713 11918 11716
rect 11860 11707 11918 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13648 11753 13676 11784
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 11146 11676 11152 11688
rect 10336 11648 11152 11676
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 13648 11676 13676 11707
rect 15010 11704 15016 11756
rect 15068 11744 15074 11756
rect 16574 11744 16580 11756
rect 15068 11716 16580 11744
rect 15068 11704 15074 11716
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17000 11716 17158 11744
rect 17000 11704 17006 11716
rect 11756 11648 13676 11676
rect 13909 11679 13967 11685
rect 11756 11636 11762 11648
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 13998 11676 14004 11688
rect 13955 11648 14004 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 16850 11676 16856 11688
rect 15703 11648 16856 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 8202 11568 8208 11620
rect 8260 11608 8266 11620
rect 8260 11580 12434 11608
rect 8260 11568 8266 11580
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6178 11540 6184 11552
rect 6043 11512 6184 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 9999 11543 10057 11549
rect 9999 11509 10011 11543
rect 10045 11540 10057 11543
rect 10410 11540 10416 11552
rect 10045 11512 10416 11540
rect 10045 11509 10057 11512
rect 9999 11503 10057 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 12406 11540 12434 11580
rect 15672 11540 15700 11639
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 18046 11636 18052 11688
rect 18104 11636 18110 11688
rect 15838 11568 15844 11620
rect 15896 11608 15902 11620
rect 17957 11611 18015 11617
rect 17957 11608 17969 11611
rect 15896 11580 17969 11608
rect 15896 11568 15902 11580
rect 17957 11577 17969 11580
rect 18003 11577 18015 11611
rect 17957 11571 18015 11577
rect 12406 11512 15700 11540
rect 18325 11543 18383 11549
rect 18325 11509 18337 11543
rect 18371 11540 18383 11543
rect 18690 11540 18696 11552
rect 18371 11512 18696 11540
rect 18371 11509 18383 11512
rect 18325 11503 18383 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 1104 11450 20700 11472
rect 1104 11398 3399 11450
rect 3451 11398 3463 11450
rect 3515 11398 3527 11450
rect 3579 11398 3591 11450
rect 3643 11398 3655 11450
rect 3707 11398 8298 11450
rect 8350 11398 8362 11450
rect 8414 11398 8426 11450
rect 8478 11398 8490 11450
rect 8542 11398 8554 11450
rect 8606 11398 13197 11450
rect 13249 11398 13261 11450
rect 13313 11398 13325 11450
rect 13377 11398 13389 11450
rect 13441 11398 13453 11450
rect 13505 11398 18096 11450
rect 18148 11398 18160 11450
rect 18212 11398 18224 11450
rect 18276 11398 18288 11450
rect 18340 11398 18352 11450
rect 18404 11398 20700 11450
rect 1104 11376 20700 11398
rect 4614 11336 4620 11348
rect 4575 11308 4620 11336
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 6822 11336 6828 11348
rect 5491 11308 6828 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 15010 11296 15016 11348
rect 15068 11336 15074 11348
rect 15197 11339 15255 11345
rect 15197 11336 15209 11339
rect 15068 11308 15209 11336
rect 15068 11296 15074 11308
rect 15197 11305 15209 11308
rect 15243 11305 15255 11339
rect 15838 11336 15844 11348
rect 15799 11308 15844 11336
rect 15197 11299 15255 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 17681 11339 17739 11345
rect 17681 11305 17693 11339
rect 17727 11336 17739 11339
rect 17770 11336 17776 11348
rect 17727 11308 17776 11336
rect 17727 11305 17739 11308
rect 17681 11299 17739 11305
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 1486 11228 1492 11280
rect 1544 11268 1550 11280
rect 1581 11271 1639 11277
rect 1581 11268 1593 11271
rect 1544 11240 1593 11268
rect 1544 11228 1550 11240
rect 1581 11237 1593 11240
rect 1627 11237 1639 11271
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 1581 11231 1639 11237
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 16853 11271 16911 11277
rect 16853 11268 16865 11271
rect 16264 11240 16865 11268
rect 16264 11228 16270 11240
rect 16853 11237 16865 11240
rect 16899 11237 16911 11271
rect 16853 11231 16911 11237
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 7929 11203 7987 11209
rect 6503 11172 7880 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 5258 11132 5264 11144
rect 5219 11104 5264 11132
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 7852 11132 7880 11172
rect 7929 11169 7941 11203
rect 7975 11200 7987 11203
rect 8110 11200 8116 11212
rect 7975 11172 8116 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 11238 11200 11244 11212
rect 10643 11172 11244 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 17954 11200 17960 11212
rect 17000 11172 17960 11200
rect 17000 11160 17006 11172
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 16028 11144 16080 11150
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 7852 11104 8585 11132
rect 8573 11101 8585 11104
rect 8619 11132 8631 11135
rect 8662 11132 8668 11144
rect 8619 11104 8668 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 11422 11141 11428 11144
rect 11400 11135 11428 11141
rect 11400 11101 11412 11135
rect 11400 11095 11428 11101
rect 11422 11092 11428 11095
rect 11480 11092 11486 11144
rect 17862 11132 17868 11144
rect 17823 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 16028 11086 16080 11092
rect 7742 11064 7748 11076
rect 7655 11036 7748 11064
rect 7742 11024 7748 11036
rect 7800 11064 7806 11076
rect 9490 11064 9496 11076
rect 7800 11036 9496 11064
rect 7800 11024 7806 11036
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 10226 11064 10232 11076
rect 9916 11036 10232 11064
rect 9916 11024 9922 11036
rect 10226 11024 10232 11036
rect 10284 11064 10290 11076
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 10284 11036 10793 11064
rect 10284 11024 10290 11036
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 10781 11027 10839 11033
rect 14921 11067 14979 11073
rect 14921 11033 14933 11067
rect 14967 11064 14979 11067
rect 15194 11064 15200 11076
rect 14967 11036 15200 11064
rect 14967 11033 14979 11036
rect 14921 11027 14979 11033
rect 15194 11024 15200 11036
rect 15252 11064 15258 11076
rect 15562 11064 15568 11076
rect 15252 11036 15568 11064
rect 15252 11024 15258 11036
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 8389 10999 8447 11005
rect 8389 10965 8401 10999
rect 8435 10996 8447 10999
rect 8662 10996 8668 11008
rect 8435 10968 8668 10996
rect 8435 10965 8447 10968
rect 8389 10959 8447 10965
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 11471 10999 11529 11005
rect 11471 10965 11483 10999
rect 11517 10996 11529 10999
rect 11882 10996 11888 11008
rect 11517 10968 11888 10996
rect 11517 10965 11529 10968
rect 11471 10959 11529 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 1104 10906 20859 10928
rect 1104 10854 5848 10906
rect 5900 10854 5912 10906
rect 5964 10854 5976 10906
rect 6028 10854 6040 10906
rect 6092 10854 6104 10906
rect 6156 10854 10747 10906
rect 10799 10854 10811 10906
rect 10863 10854 10875 10906
rect 10927 10854 10939 10906
rect 10991 10854 11003 10906
rect 11055 10854 15646 10906
rect 15698 10854 15710 10906
rect 15762 10854 15774 10906
rect 15826 10854 15838 10906
rect 15890 10854 15902 10906
rect 15954 10854 20545 10906
rect 20597 10854 20609 10906
rect 20661 10854 20673 10906
rect 20725 10854 20737 10906
rect 20789 10854 20801 10906
rect 20853 10854 20859 10906
rect 1104 10832 20859 10854
rect 3970 10792 3976 10804
rect 3931 10764 3976 10792
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 17957 10795 18015 10801
rect 17957 10792 17969 10795
rect 17920 10764 17969 10792
rect 17920 10752 17926 10764
rect 17957 10761 17969 10764
rect 18003 10761 18015 10795
rect 17957 10755 18015 10761
rect 8754 10724 8760 10736
rect 8588 10696 8760 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2314 10656 2320 10668
rect 2271 10628 2320 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3292 10628 3341 10656
rect 3292 10616 3298 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10656 7803 10659
rect 8202 10656 8208 10668
rect 7791 10628 8208 10656
rect 7791 10625 7803 10628
rect 7745 10619 7803 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8588 10665 8616 10696
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 10781 10727 10839 10733
rect 10781 10724 10793 10727
rect 10074 10710 10793 10724
rect 10060 10696 10793 10710
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7432 10560 7665 10588
rect 7432 10548 7438 10560
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 7653 10551 7711 10557
rect 8680 10560 8861 10588
rect 8113 10523 8171 10529
rect 8113 10489 8125 10523
rect 8159 10520 8171 10523
rect 8680 10520 8708 10560
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 10060 10588 10088 10696
rect 10781 10693 10793 10696
rect 10827 10693 10839 10727
rect 10781 10687 10839 10693
rect 12618 10684 12624 10736
rect 12676 10684 12682 10736
rect 14642 10684 14648 10736
rect 14700 10684 14706 10736
rect 18690 10724 18696 10736
rect 18651 10696 18696 10724
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 19334 10684 19340 10736
rect 19392 10684 19398 10736
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11606 10656 11612 10668
rect 11011 10628 11612 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 13906 10656 13912 10668
rect 13867 10628 13912 10656
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 17770 10656 17776 10668
rect 17731 10628 17776 10656
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 11698 10588 11704 10600
rect 9272 10560 10088 10588
rect 11659 10560 11704 10588
rect 9272 10548 9278 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 11974 10588 11980 10600
rect 11935 10560 11980 10588
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10588 18478 10600
rect 18782 10588 18788 10600
rect 18472 10560 18788 10588
rect 18472 10548 18478 10560
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 8159 10492 8708 10520
rect 8159 10489 8171 10492
rect 8113 10483 8171 10489
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 1946 10452 1952 10464
rect 1811 10424 1952 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2832 10424 2881 10452
rect 2832 10412 2838 10424
rect 2869 10421 2881 10424
rect 2915 10421 2927 10455
rect 2869 10415 2927 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9640 10424 10333 10452
rect 9640 10412 9646 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 13449 10455 13507 10461
rect 13449 10421 13461 10455
rect 13495 10452 13507 10455
rect 14274 10452 14280 10464
rect 13495 10424 14280 10452
rect 13495 10421 13507 10424
rect 13449 10415 13507 10421
rect 14274 10412 14280 10424
rect 14332 10412 14338 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 15620 10424 15669 10452
rect 15620 10412 15626 10424
rect 15657 10421 15669 10424
rect 15703 10421 15715 10455
rect 20162 10452 20168 10464
rect 20123 10424 20168 10452
rect 15657 10415 15715 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 1104 10362 20700 10384
rect 1104 10310 3399 10362
rect 3451 10310 3463 10362
rect 3515 10310 3527 10362
rect 3579 10310 3591 10362
rect 3643 10310 3655 10362
rect 3707 10310 8298 10362
rect 8350 10310 8362 10362
rect 8414 10310 8426 10362
rect 8478 10310 8490 10362
rect 8542 10310 8554 10362
rect 8606 10310 13197 10362
rect 13249 10310 13261 10362
rect 13313 10310 13325 10362
rect 13377 10310 13389 10362
rect 13441 10310 13453 10362
rect 13505 10310 18096 10362
rect 18148 10310 18160 10362
rect 18212 10310 18224 10362
rect 18276 10310 18288 10362
rect 18340 10310 18352 10362
rect 18404 10310 20700 10362
rect 1104 10288 20700 10310
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3292 10220 3433 10248
rect 3292 10208 3298 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 11422 10248 11428 10260
rect 11383 10220 11428 10248
rect 3421 10211 3479 10217
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 12253 10251 12311 10257
rect 12253 10217 12265 10251
rect 12299 10248 12311 10251
rect 12618 10248 12624 10260
rect 12299 10220 12624 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 16022 10248 16028 10260
rect 15983 10220 16028 10248
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 11882 10180 11888 10192
rect 11843 10152 11888 10180
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 11057 10115 11115 10121
rect 11057 10112 11069 10115
rect 9600 10084 11069 10112
rect 9600 10056 9628 10084
rect 11057 10081 11069 10084
rect 11103 10081 11115 10115
rect 11057 10075 11115 10081
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11664 10084 12081 10112
rect 11664 10072 11670 10084
rect 12069 10081 12081 10084
rect 12115 10112 12127 10115
rect 15194 10112 15200 10124
rect 12115 10084 15200 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 8113 10047 8171 10053
rect 2832 10016 2877 10044
rect 2832 10004 2838 10016
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8662 10044 8668 10056
rect 8159 10016 8668 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9376 10047 9434 10053
rect 9376 10013 9388 10047
rect 9422 10044 9434 10047
rect 9582 10044 9588 10056
rect 9422 10016 9588 10044
rect 9422 10013 9434 10016
rect 9376 10007 9434 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9950 10044 9956 10056
rect 9911 10016 9956 10044
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10594 10044 10600 10056
rect 10507 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10044 10658 10056
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 10652 10016 11253 10044
rect 10652 10004 10658 10016
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 11241 10007 11299 10013
rect 12406 10016 14289 10044
rect 12406 9976 12434 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 20162 10044 20168 10056
rect 20123 10016 20168 10044
rect 14277 10007 14335 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 14550 9976 14556 9988
rect 9324 9948 12434 9976
rect 14463 9948 14556 9976
rect 9324 9920 9352 9948
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 15194 9936 15200 9988
rect 15252 9936 15258 9988
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8754 9908 8760 9920
rect 8343 9880 8760 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8754 9868 8760 9880
rect 8812 9908 8818 9920
rect 9306 9908 9312 9920
rect 8812 9880 9312 9908
rect 8812 9868 8818 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9447 9911 9505 9917
rect 9447 9877 9459 9911
rect 9493 9908 9505 9911
rect 10502 9908 10508 9920
rect 9493 9880 10508 9908
rect 9493 9877 9505 9880
rect 9447 9871 9505 9877
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 14568 9908 14596 9936
rect 12032 9880 14596 9908
rect 12032 9868 12038 9880
rect 1104 9818 20859 9840
rect 1104 9766 5848 9818
rect 5900 9766 5912 9818
rect 5964 9766 5976 9818
rect 6028 9766 6040 9818
rect 6092 9766 6104 9818
rect 6156 9766 10747 9818
rect 10799 9766 10811 9818
rect 10863 9766 10875 9818
rect 10927 9766 10939 9818
rect 10991 9766 11003 9818
rect 11055 9766 15646 9818
rect 15698 9766 15710 9818
rect 15762 9766 15774 9818
rect 15826 9766 15838 9818
rect 15890 9766 15902 9818
rect 15954 9766 20545 9818
rect 20597 9766 20609 9818
rect 20661 9766 20673 9818
rect 20725 9766 20737 9818
rect 20789 9766 20801 9818
rect 20853 9766 20859 9818
rect 1104 9744 20859 9766
rect 9950 9704 9956 9716
rect 9911 9676 9956 9704
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 17770 9704 17776 9716
rect 17731 9676 17776 9704
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 4755 9639 4813 9645
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 2041 9571 2099 9577
rect 2041 9568 2053 9571
rect 1912 9540 2053 9568
rect 1912 9528 1918 9540
rect 2041 9537 2053 9540
rect 2087 9537 2099 9571
rect 4356 9568 4384 9622
rect 4755 9605 4767 9639
rect 4801 9636 4813 9639
rect 4890 9636 4896 9648
rect 4801 9608 4896 9636
rect 4801 9605 4813 9608
rect 4755 9599 4813 9605
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 10560 9608 10732 9636
rect 10560 9596 10566 9608
rect 5534 9568 5540 9580
rect 4356 9540 5540 9568
rect 2041 9531 2099 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 10594 9568 10600 9580
rect 10555 9540 10600 9568
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10704 9577 10732 9608
rect 17218 9596 17224 9648
rect 17276 9636 17282 9648
rect 18693 9639 18751 9645
rect 18693 9636 18705 9639
rect 17276 9608 18705 9636
rect 17276 9596 17282 9608
rect 18693 9605 18705 9608
rect 18739 9605 18751 9639
rect 18693 9599 18751 9605
rect 19334 9596 19340 9648
rect 19392 9596 19398 9648
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 17954 9568 17960 9580
rect 17915 9540 17960 9568
rect 10689 9531 10747 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 1670 9500 1676 9512
rect 1631 9472 1676 9500
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 3292 9472 3341 9500
rect 3292 9460 3298 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 11974 9500 11980 9512
rect 4580 9472 11980 9500
rect 4580 9460 4586 9472
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18414 9500 18420 9512
rect 17920 9472 18420 9500
rect 17920 9460 17926 9472
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 7282 9364 7288 9376
rect 6963 9336 7288 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 10410 9364 10416 9376
rect 10371 9336 10416 9364
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 1104 9274 20700 9296
rect 1104 9222 3399 9274
rect 3451 9222 3463 9274
rect 3515 9222 3527 9274
rect 3579 9222 3591 9274
rect 3643 9222 3655 9274
rect 3707 9222 8298 9274
rect 8350 9222 8362 9274
rect 8414 9222 8426 9274
rect 8478 9222 8490 9274
rect 8542 9222 8554 9274
rect 8606 9222 13197 9274
rect 13249 9222 13261 9274
rect 13313 9222 13325 9274
rect 13377 9222 13389 9274
rect 13441 9222 13453 9274
rect 13505 9222 18096 9274
rect 18148 9222 18160 9274
rect 18212 9222 18224 9274
rect 18276 9222 18288 9274
rect 18340 9222 18352 9274
rect 18404 9222 20700 9274
rect 1104 9200 20700 9222
rect 3234 9120 3240 9172
rect 3292 9169 3298 9172
rect 3292 9163 3341 9169
rect 3292 9129 3295 9163
rect 3329 9129 3341 9163
rect 3292 9123 3341 9129
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7466 9160 7472 9172
rect 6871 9132 7472 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 3292 9120 3298 9123
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 18012 9132 18061 9160
rect 18012 9120 18018 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 12713 9095 12771 9101
rect 12713 9061 12725 9095
rect 12759 9092 12771 9095
rect 13814 9092 13820 9104
rect 12759 9064 13820 9092
rect 12759 9061 12771 9064
rect 12713 9055 12771 9061
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 19429 9095 19487 9101
rect 19429 9092 19441 9095
rect 17920 9064 19441 9092
rect 17920 9052 17926 9064
rect 19429 9061 19441 9064
rect 19475 9061 19487 9095
rect 19429 9055 19487 9061
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 9582 9024 9588 9036
rect 3200 8996 9588 9024
rect 3200 8984 3206 8996
rect 9582 8984 9588 8996
rect 9640 9024 9646 9036
rect 12250 9024 12256 9036
rect 9640 8996 12256 9024
rect 9640 8984 9646 8996
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 9024 15439 9027
rect 16022 9024 16028 9036
rect 15427 8996 16028 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16853 9027 16911 9033
rect 16853 8993 16865 9027
rect 16899 8993 16911 9027
rect 16853 8987 16911 8993
rect 3386 8959 3444 8965
rect 3386 8925 3398 8959
rect 3432 8956 3444 8959
rect 4522 8956 4528 8968
rect 3432 8928 4384 8956
rect 4483 8928 4528 8956
rect 3432 8925 3444 8928
rect 3386 8919 3444 8925
rect 4356 8832 4384 8928
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 7282 8956 7288 8968
rect 7195 8928 7288 8956
rect 5077 8919 5135 8925
rect 5092 8888 5120 8919
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 8110 8956 8116 8968
rect 8071 8928 8116 8956
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10318 8956 10324 8968
rect 9907 8928 10324 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 12066 8916 12072 8968
rect 12124 8956 12130 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12124 8928 12541 8956
rect 12124 8916 12130 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 13538 8956 13544 8968
rect 13495 8928 13544 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 15102 8956 15108 8968
rect 15063 8928 15108 8956
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 16868 8956 16896 8987
rect 17126 8956 17132 8968
rect 16868 8928 17132 8956
rect 17126 8916 17132 8928
rect 17184 8956 17190 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 17184 8928 17325 8956
rect 17184 8916 17190 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18414 8956 18420 8968
rect 18375 8928 18420 8956
rect 18233 8919 18291 8925
rect 5258 8888 5264 8900
rect 5092 8860 5264 8888
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5442 8888 5448 8900
rect 5399 8860 5448 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 6914 8888 6920 8900
rect 6578 8860 6920 8888
rect 6914 8848 6920 8860
rect 6972 8848 6978 8900
rect 7300 8888 7328 8916
rect 9950 8888 9956 8900
rect 7300 8860 9956 8888
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 17586 8888 17592 8900
rect 16606 8860 17592 8888
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 7466 8820 7472 8832
rect 7427 8792 7472 8820
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7926 8820 7932 8832
rect 7887 8792 7932 8820
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9766 8820 9772 8832
rect 9723 8792 9772 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 12860 8792 13277 8820
rect 12860 8780 12866 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16684 8820 16712 8860
rect 17586 8848 17592 8860
rect 17644 8848 17650 8900
rect 18248 8888 18276 8919
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 19334 8888 19340 8900
rect 18248 8860 19340 8888
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 19610 8888 19616 8900
rect 19571 8860 19616 8888
rect 19610 8848 19616 8860
rect 19668 8848 19674 8900
rect 16172 8792 16712 8820
rect 17497 8823 17555 8829
rect 16172 8780 16178 8792
rect 17497 8789 17509 8823
rect 17543 8820 17555 8823
rect 19242 8820 19248 8832
rect 17543 8792 19248 8820
rect 17543 8789 17555 8792
rect 17497 8783 17555 8789
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 1104 8730 20859 8752
rect 1104 8678 5848 8730
rect 5900 8678 5912 8730
rect 5964 8678 5976 8730
rect 6028 8678 6040 8730
rect 6092 8678 6104 8730
rect 6156 8678 10747 8730
rect 10799 8678 10811 8730
rect 10863 8678 10875 8730
rect 10927 8678 10939 8730
rect 10991 8678 11003 8730
rect 11055 8678 15646 8730
rect 15698 8678 15710 8730
rect 15762 8678 15774 8730
rect 15826 8678 15838 8730
rect 15890 8678 15902 8730
rect 15954 8678 20545 8730
rect 20597 8678 20609 8730
rect 20661 8678 20673 8730
rect 20725 8678 20737 8730
rect 20789 8678 20801 8730
rect 20853 8678 20859 8730
rect 1104 8656 20859 8678
rect 2498 8616 2504 8628
rect 2459 8588 2504 8616
rect 2498 8576 2504 8588
rect 2556 8616 2562 8628
rect 2774 8616 2780 8628
rect 2556 8588 2780 8616
rect 2556 8576 2562 8588
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 5258 8616 5264 8628
rect 4080 8588 5264 8616
rect 4080 8548 4108 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5718 8616 5724 8628
rect 5679 8588 5724 8616
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 12066 8616 12072 8628
rect 12027 8588 12072 8616
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 15381 8619 15439 8625
rect 15381 8616 15393 8619
rect 15160 8588 15393 8616
rect 15160 8576 15166 8588
rect 15381 8585 15393 8588
rect 15427 8585 15439 8619
rect 19978 8616 19984 8628
rect 19939 8588 19984 8616
rect 15381 8579 15439 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 3988 8520 4108 8548
rect 3988 8489 4016 8520
rect 4798 8508 4804 8560
rect 4856 8508 4862 8560
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 7926 8548 7932 8560
rect 6779 8520 7932 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 7926 8508 7932 8520
rect 7984 8508 7990 8560
rect 8389 8551 8447 8557
rect 8389 8517 8401 8551
rect 8435 8548 8447 8551
rect 8662 8548 8668 8560
rect 8435 8520 8668 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 12802 8548 12808 8560
rect 12544 8520 12808 8548
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 3973 8443 4031 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 10318 8480 10324 8492
rect 10279 8452 10324 8480
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 12544 8489 12572 8520
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 15654 8548 15660 8560
rect 14030 8520 15660 8548
rect 15654 8508 15660 8520
rect 15712 8548 15718 8560
rect 16114 8548 16120 8560
rect 15712 8520 16120 8548
rect 15712 8508 15718 8520
rect 16114 8508 16120 8520
rect 16172 8508 16178 8560
rect 17126 8548 17132 8560
rect 17087 8520 17132 8548
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17586 8508 17592 8560
rect 17644 8508 17650 8560
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12529 8483 12587 8489
rect 11931 8452 12434 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12406 8424 12434 8452
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 15565 8483 15623 8489
rect 15565 8480 15577 8483
rect 14737 8443 14795 8449
rect 14936 8452 15577 8480
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 3142 8412 3148 8424
rect 2731 8384 3148 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 4246 8412 4252 8424
rect 4207 8384 4252 8412
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8381 8171 8415
rect 12406 8384 12440 8424
rect 8113 8375 8171 8381
rect 2866 8344 2872 8356
rect 2827 8316 2872 8344
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 5408 8316 6561 8344
rect 5408 8304 5414 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 7653 8347 7711 8353
rect 7653 8313 7665 8347
rect 7699 8344 7711 8347
rect 8128 8344 8156 8375
rect 12434 8372 12440 8384
rect 12492 8412 12498 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12492 8384 12817 8412
rect 12492 8372 12498 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 14752 8412 14780 8443
rect 12952 8384 14780 8412
rect 12952 8372 12958 8384
rect 14936 8353 14964 8452
rect 15565 8449 15577 8452
rect 15611 8480 15623 8483
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 15611 8452 16037 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 16025 8449 16037 8452
rect 16071 8449 16083 8483
rect 19242 8480 19248 8492
rect 19203 8452 19248 8480
rect 16025 8443 16083 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 20162 8480 20168 8492
rect 20123 8452 20168 8480
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 7699 8316 8156 8344
rect 14921 8347 14979 8353
rect 7699 8313 7711 8316
rect 7653 8307 7711 8313
rect 14921 8313 14933 8347
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 16868 8344 16896 8375
rect 16255 8316 16896 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9861 8279 9919 8285
rect 9861 8276 9873 8279
rect 9732 8248 9873 8276
rect 9732 8236 9738 8248
rect 9861 8245 9873 8248
rect 9907 8245 9919 8279
rect 10502 8276 10508 8288
rect 10463 8248 10508 8276
rect 9861 8239 9919 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 14277 8279 14335 8285
rect 14277 8245 14289 8279
rect 14323 8276 14335 8279
rect 14550 8276 14556 8288
rect 14323 8248 14556 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 17770 8236 17776 8288
rect 17828 8276 17834 8288
rect 18601 8279 18659 8285
rect 18601 8276 18613 8279
rect 17828 8248 18613 8276
rect 17828 8236 17834 8248
rect 18601 8245 18613 8248
rect 18647 8245 18659 8279
rect 19058 8276 19064 8288
rect 19019 8248 19064 8276
rect 18601 8239 18659 8245
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 1104 8186 20700 8208
rect 1104 8134 3399 8186
rect 3451 8134 3463 8186
rect 3515 8134 3527 8186
rect 3579 8134 3591 8186
rect 3643 8134 3655 8186
rect 3707 8134 8298 8186
rect 8350 8134 8362 8186
rect 8414 8134 8426 8186
rect 8478 8134 8490 8186
rect 8542 8134 8554 8186
rect 8606 8134 13197 8186
rect 13249 8134 13261 8186
rect 13313 8134 13325 8186
rect 13377 8134 13389 8186
rect 13441 8134 13453 8186
rect 13505 8134 18096 8186
rect 18148 8134 18160 8186
rect 18212 8134 18224 8186
rect 18276 8134 18288 8186
rect 18340 8134 18352 8186
rect 18404 8134 20700 8186
rect 1104 8112 20700 8134
rect 4246 8081 4252 8084
rect 4203 8075 4252 8081
rect 4203 8041 4215 8075
rect 4249 8041 4252 8075
rect 4203 8035 4252 8041
rect 4246 8032 4252 8035
rect 4304 8032 4310 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 8573 8075 8631 8081
rect 7616 8044 8524 8072
rect 7616 8032 7622 8044
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 3234 8004 3240 8016
rect 3099 7976 3240 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3234 7964 3240 7976
rect 3292 7964 3298 8016
rect 5307 7939 5365 7945
rect 5307 7905 5319 7939
rect 5353 7936 5365 7939
rect 5442 7936 5448 7948
rect 5353 7908 5448 7936
rect 5353 7905 5365 7908
rect 5307 7899 5365 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 8110 7936 8116 7948
rect 7147 7908 8116 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8496 7936 8524 8044
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8662 8072 8668 8084
rect 8619 8044 8668 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 10318 8072 10324 8084
rect 9907 8044 10324 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 10952 8075 11010 8081
rect 10952 8041 10964 8075
rect 10998 8072 11010 8075
rect 11146 8072 11152 8084
rect 10998 8044 11152 8072
rect 10998 8041 11010 8044
rect 10952 8035 11010 8041
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 13081 8075 13139 8081
rect 12492 8044 12537 8072
rect 12492 8032 12498 8044
rect 13081 8041 13093 8075
rect 13127 8072 13139 8075
rect 13538 8072 13544 8084
rect 13127 8044 13544 8072
rect 13127 8041 13139 8044
rect 13081 8035 13139 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 16022 8072 16028 8084
rect 15983 8044 16028 8072
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 17313 8075 17371 8081
rect 17313 8041 17325 8075
rect 17359 8072 17371 8075
rect 18506 8072 18512 8084
rect 17359 8044 18512 8072
rect 17359 8041 17371 8044
rect 17313 8035 17371 8041
rect 18506 8032 18512 8044
rect 18564 8072 18570 8084
rect 19610 8072 19616 8084
rect 18564 8044 19616 8072
rect 18564 8032 18570 8044
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 9950 8004 9956 8016
rect 9692 7976 9956 8004
rect 8496 7908 9628 7936
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1728 7840 1777 7868
rect 1728 7828 1734 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 3142 7828 3148 7880
rect 3200 7868 3206 7880
rect 4338 7877 4344 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 3200 7840 3249 7868
rect 3200 7828 3206 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 4306 7871 4344 7877
rect 4306 7868 4318 7871
rect 4251 7840 4318 7868
rect 3237 7831 3295 7837
rect 4306 7837 4318 7840
rect 4396 7868 4402 7880
rect 5220 7871 5278 7877
rect 5220 7868 5232 7871
rect 4396 7840 5232 7868
rect 4306 7831 4344 7837
rect 4338 7828 4344 7831
rect 4396 7828 4402 7840
rect 5220 7837 5232 7840
rect 5266 7868 5278 7871
rect 5626 7868 5632 7880
rect 5266 7840 5632 7868
rect 5266 7837 5278 7840
rect 5220 7831 5278 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 6822 7868 6828 7880
rect 6783 7840 6828 7868
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 9490 7800 9496 7812
rect 8326 7772 9496 7800
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 9600 7800 9628 7908
rect 9692 7877 9720 7976
rect 9950 7964 9956 7976
rect 10008 8004 10014 8016
rect 13725 8007 13783 8013
rect 10008 7976 10824 8004
rect 10008 7964 10014 7976
rect 10502 7896 10508 7948
rect 10560 7936 10566 7948
rect 10689 7939 10747 7945
rect 10689 7936 10701 7939
rect 10560 7908 10701 7936
rect 10560 7896 10566 7908
rect 10689 7905 10701 7908
rect 10735 7905 10747 7939
rect 10796 7936 10824 7976
rect 13725 7973 13737 8007
rect 13771 8004 13783 8007
rect 16669 8007 16727 8013
rect 13771 7976 14320 8004
rect 13771 7973 13783 7976
rect 13725 7967 13783 7973
rect 14292 7945 14320 7976
rect 16669 7973 16681 8007
rect 16715 7973 16727 8007
rect 18414 8004 18420 8016
rect 18375 7976 18420 8004
rect 16669 7967 16727 7973
rect 14277 7939 14335 7945
rect 10796 7908 12434 7936
rect 10689 7899 10747 7905
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 12406 7868 12434 7908
rect 14277 7905 14289 7939
rect 14323 7905 14335 7939
rect 14550 7936 14556 7948
rect 14511 7908 14556 7936
rect 14277 7899 14335 7905
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 12894 7868 12900 7880
rect 12406 7840 12900 7868
rect 9677 7831 9735 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 15654 7828 15660 7880
rect 15712 7828 15718 7880
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 16080 7840 16497 7868
rect 16080 7828 16086 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16684 7868 16712 7967
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 19429 8007 19487 8013
rect 19429 7973 19441 8007
rect 19475 7973 19487 8007
rect 19429 7967 19487 7973
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7936 18199 7939
rect 19444 7936 19472 7967
rect 18187 7908 19472 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 17129 7871 17187 7877
rect 17129 7868 17141 7871
rect 16684 7840 17141 7868
rect 16485 7831 16543 7837
rect 17129 7837 17141 7840
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 19058 7868 19064 7880
rect 18095 7840 19064 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19610 7868 19616 7880
rect 19571 7840 19616 7868
rect 19610 7828 19616 7840
rect 19668 7828 19674 7880
rect 9600 7772 11454 7800
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2409 7735 2467 7741
rect 2409 7732 2421 7735
rect 2372 7704 2421 7732
rect 2372 7692 2378 7704
rect 2409 7701 2421 7704
rect 2455 7701 2467 7735
rect 2409 7695 2467 7701
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3970 7732 3976 7744
rect 3467 7704 3976 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 11348 7732 11376 7772
rect 15672 7732 15700 7828
rect 11348 7704 15700 7732
rect 1104 7642 20859 7664
rect 1104 7590 5848 7642
rect 5900 7590 5912 7642
rect 5964 7590 5976 7642
rect 6028 7590 6040 7642
rect 6092 7590 6104 7642
rect 6156 7590 10747 7642
rect 10799 7590 10811 7642
rect 10863 7590 10875 7642
rect 10927 7590 10939 7642
rect 10991 7590 11003 7642
rect 11055 7590 15646 7642
rect 15698 7590 15710 7642
rect 15762 7590 15774 7642
rect 15826 7590 15838 7642
rect 15890 7590 15902 7642
rect 15954 7590 20545 7642
rect 20597 7590 20609 7642
rect 20661 7590 20673 7642
rect 20725 7590 20737 7642
rect 20789 7590 20801 7642
rect 20853 7590 20859 7642
rect 1104 7568 20859 7590
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 7193 7531 7251 7537
rect 7193 7528 7205 7531
rect 6880 7500 7205 7528
rect 6880 7488 6886 7500
rect 7193 7497 7205 7500
rect 7239 7497 7251 7531
rect 7193 7491 7251 7497
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 11146 7528 11152 7540
rect 9548 7500 9812 7528
rect 11107 7500 11152 7528
rect 9548 7488 9554 7500
rect 2498 7420 2504 7472
rect 2556 7420 2562 7472
rect 9674 7460 9680 7472
rect 9635 7432 9680 7460
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 9784 7460 9812 7500
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 17957 7531 18015 7537
rect 17957 7497 17969 7531
rect 18003 7528 18015 7531
rect 19610 7528 19616 7540
rect 18003 7500 19616 7528
rect 18003 7497 18015 7500
rect 17957 7491 18015 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 9784 7432 10166 7460
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5684 7364 6009 7392
rect 5684 7352 5690 7364
rect 5997 7361 6009 7364
rect 6043 7392 6055 7395
rect 7282 7392 7288 7404
rect 6043 7364 7288 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7466 7392 7472 7404
rect 7423 7364 7472 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8662 7392 8668 7404
rect 8619 7364 8668 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 11164 7392 11192 7488
rect 19334 7420 19340 7472
rect 19392 7420 19398 7472
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11164 7364 11897 7392
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14608 7364 14841 7392
rect 14608 7352 14614 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 17770 7392 17776 7404
rect 17731 7364 17776 7392
rect 14829 7355 14887 7361
rect 17770 7352 17776 7364
rect 17828 7352 17834 7404
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 1854 7324 1860 7336
rect 1627 7296 1716 7324
rect 1815 7296 1860 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 1688 7200 1716 7296
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 5534 7324 5540 7336
rect 4571 7296 5540 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 5534 7284 5540 7296
rect 5592 7324 5598 7336
rect 5718 7324 5724 7336
rect 5592 7296 5724 7324
rect 5592 7284 5598 7296
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 9766 7324 9772 7336
rect 9447 7296 9772 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 17126 7284 17132 7336
rect 17184 7324 17190 7336
rect 17862 7324 17868 7336
rect 17184 7296 17868 7324
rect 17184 7284 17190 7296
rect 17862 7284 17868 7296
rect 17920 7324 17926 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 17920 7296 18429 7324
rect 17920 7284 17926 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18690 7324 18696 7336
rect 18651 7296 18696 7324
rect 18417 7287 18475 7293
rect 18690 7284 18696 7296
rect 18748 7284 18754 7336
rect 4338 7256 4344 7268
rect 4299 7228 4344 7256
rect 4338 7216 4344 7228
rect 4396 7216 4402 7268
rect 4448 7228 5672 7256
rect 1670 7148 1676 7200
rect 1728 7148 1734 7200
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 3292 7160 3341 7188
rect 3292 7148 3298 7160
rect 3329 7157 3341 7160
rect 3375 7157 3387 7191
rect 3329 7151 3387 7157
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4448 7188 4476 7228
rect 5644 7200 5672 7228
rect 3844 7160 4476 7188
rect 4709 7191 4767 7197
rect 3844 7148 3850 7160
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4798 7188 4804 7200
rect 4755 7160 4804 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5684 7160 5825 7188
rect 5684 7148 5690 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 8757 7191 8815 7197
rect 8757 7157 8769 7191
rect 8803 7188 8815 7191
rect 9122 7188 9128 7200
rect 8803 7160 9128 7188
rect 8803 7157 8815 7160
rect 8757 7151 8815 7157
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 11480 7160 11713 7188
rect 11480 7148 11486 7160
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 15013 7191 15071 7197
rect 15013 7157 15025 7191
rect 15059 7188 15071 7191
rect 15654 7188 15660 7200
rect 15059 7160 15660 7188
rect 15059 7157 15071 7160
rect 15013 7151 15071 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 20162 7188 20168 7200
rect 20123 7160 20168 7188
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 1104 7098 20700 7120
rect 1104 7046 3399 7098
rect 3451 7046 3463 7098
rect 3515 7046 3527 7098
rect 3579 7046 3591 7098
rect 3643 7046 3655 7098
rect 3707 7046 8298 7098
rect 8350 7046 8362 7098
rect 8414 7046 8426 7098
rect 8478 7046 8490 7098
rect 8542 7046 8554 7098
rect 8606 7046 13197 7098
rect 13249 7046 13261 7098
rect 13313 7046 13325 7098
rect 13377 7046 13389 7098
rect 13441 7046 13453 7098
rect 13505 7046 18096 7098
rect 18148 7046 18160 7098
rect 18212 7046 18224 7098
rect 18276 7046 18288 7098
rect 18340 7046 18352 7098
rect 18404 7046 20700 7098
rect 1104 7024 20700 7046
rect 2961 6987 3019 6993
rect 2961 6953 2973 6987
rect 3007 6984 3019 6987
rect 3142 6984 3148 6996
rect 3007 6956 3148 6984
rect 3007 6953 3019 6956
rect 2961 6947 3019 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 4111 6987 4169 6993
rect 4111 6953 4123 6987
rect 4157 6984 4169 6987
rect 4338 6984 4344 6996
rect 4157 6956 4344 6984
rect 4157 6953 4169 6956
rect 4111 6947 4169 6953
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 11241 6987 11299 6993
rect 11241 6984 11253 6987
rect 5460 6956 11253 6984
rect 1670 6876 1676 6928
rect 1728 6916 1734 6928
rect 5460 6916 5488 6956
rect 11241 6953 11253 6956
rect 11287 6984 11299 6987
rect 12342 6984 12348 6996
rect 11287 6956 12348 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 1728 6888 5488 6916
rect 1728 6876 1734 6888
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 13814 6916 13820 6928
rect 12308 6888 13820 6916
rect 12308 6876 12314 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 9214 6848 9220 6860
rect 5776 6820 9220 6848
rect 5776 6808 5782 6820
rect 2314 6780 2320 6792
rect 2275 6752 2320 6780
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3970 6740 3976 6792
rect 4028 6789 4034 6792
rect 4028 6783 4066 6789
rect 4054 6749 4066 6783
rect 5350 6780 5356 6792
rect 5311 6752 5356 6780
rect 4028 6743 4066 6749
rect 4028 6740 4034 6743
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 6748 6766 6776 6820
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9122 6780 9128 6792
rect 9083 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9732 6752 9873 6780
rect 9732 6740 9738 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 11422 6780 11428 6792
rect 11383 6752 11428 6780
rect 9861 6743 9919 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 20162 6780 20168 6792
rect 20123 6752 20168 6780
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 7377 6715 7435 6721
rect 7377 6681 7389 6715
rect 7423 6712 7435 6715
rect 7466 6712 7472 6724
rect 7423 6684 7472 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 7466 6672 7472 6684
rect 7524 6712 7530 6724
rect 15286 6712 15292 6724
rect 7524 6684 15292 6712
rect 7524 6672 7530 6684
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 7984 6616 9321 6644
rect 7984 6604 7990 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9309 6607 9367 6613
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10594 6644 10600 6656
rect 10091 6616 10600 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6644 15899 6647
rect 16850 6644 16856 6656
rect 15887 6616 16856 6644
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 1104 6554 20859 6576
rect 1104 6502 5848 6554
rect 5900 6502 5912 6554
rect 5964 6502 5976 6554
rect 6028 6502 6040 6554
rect 6092 6502 6104 6554
rect 6156 6502 10747 6554
rect 10799 6502 10811 6554
rect 10863 6502 10875 6554
rect 10927 6502 10939 6554
rect 10991 6502 11003 6554
rect 11055 6502 15646 6554
rect 15698 6502 15710 6554
rect 15762 6502 15774 6554
rect 15826 6502 15838 6554
rect 15890 6502 15902 6554
rect 15954 6502 20545 6554
rect 20597 6502 20609 6554
rect 20661 6502 20673 6554
rect 20725 6502 20737 6554
rect 20789 6502 20801 6554
rect 20853 6502 20859 6554
rect 1104 6480 20859 6502
rect 2866 6400 2872 6452
rect 2924 6449 2930 6452
rect 2924 6443 2973 6449
rect 2924 6409 2927 6443
rect 2961 6409 2973 6443
rect 7466 6440 7472 6452
rect 2924 6403 2973 6409
rect 3804 6412 7472 6440
rect 2924 6400 2930 6403
rect 3804 6372 3832 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 14093 6443 14151 6449
rect 14093 6409 14105 6443
rect 14139 6440 14151 6443
rect 15378 6440 15384 6452
rect 14139 6412 15384 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 16301 6443 16359 6449
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 18690 6440 18696 6452
rect 16347 6412 18696 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 10502 6372 10508 6384
rect 2240 6344 3832 6372
rect 3896 6344 10508 6372
rect 2240 6313 2268 6344
rect 2884 6316 2912 6344
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2866 6264 2872 6316
rect 2924 6264 2930 6316
rect 3018 6307 3076 6313
rect 3018 6273 3030 6307
rect 3064 6304 3076 6307
rect 3234 6304 3240 6316
rect 3064 6276 3240 6304
rect 3064 6273 3076 6276
rect 3018 6267 3076 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3896 6313 3924 6344
rect 10502 6332 10508 6344
rect 10560 6332 10566 6384
rect 12526 6332 12532 6384
rect 12584 6372 12590 6384
rect 12584 6344 13110 6372
rect 12584 6332 12590 6344
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 17034 6372 17040 6384
rect 16632 6344 17040 6372
rect 16632 6332 16638 6344
rect 17034 6332 17040 6344
rect 17092 6372 17098 6384
rect 17092 6344 17618 6372
rect 17092 6332 17098 6344
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 3970 6304 3976 6316
rect 3927 6276 3976 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 9214 6304 9220 6316
rect 9175 6276 9220 6304
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 10594 6304 10600 6316
rect 10555 6276 10600 6304
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 12342 6304 12348 6316
rect 12303 6276 12348 6304
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 16850 6304 16856 6316
rect 13964 6276 15134 6304
rect 16811 6276 16856 6304
rect 13964 6264 13970 6276
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 3142 6236 3148 6248
rect 2363 6208 3148 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 3142 6196 3148 6208
rect 3200 6236 3206 6248
rect 3786 6236 3792 6248
rect 3200 6208 3792 6236
rect 3200 6196 3206 6208
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 5258 6236 5264 6248
rect 5219 6208 5264 6236
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 9950 6236 9956 6248
rect 9911 6208 9956 6236
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 14182 6236 14188 6248
rect 12667 6208 14188 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 17129 6239 17187 6245
rect 17129 6236 17141 6239
rect 16132 6208 17141 6236
rect 16132 6180 16160 6208
rect 17129 6205 17141 6208
rect 17175 6205 17187 6239
rect 17129 6199 17187 6205
rect 5074 6168 5080 6180
rect 5035 6140 5080 6168
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 9766 6168 9772 6180
rect 9727 6140 9772 6168
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 15010 6128 15016 6180
rect 15068 6168 15074 6180
rect 15933 6171 15991 6177
rect 15933 6168 15945 6171
rect 15068 6140 15945 6168
rect 15068 6128 15074 6140
rect 15933 6137 15945 6140
rect 15979 6137 15991 6171
rect 15933 6131 15991 6137
rect 16114 6128 16120 6180
rect 16172 6128 16178 6180
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5626 6100 5632 6112
rect 5491 6072 5632 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8812 6072 8953 6100
rect 8812 6060 8818 6072
rect 8941 6069 8953 6072
rect 8987 6069 8999 6103
rect 8941 6063 8999 6069
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9732 6072 10149 6100
rect 9732 6060 9738 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10560 6072 10793 6100
rect 10560 6060 10566 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 10781 6063 10839 6069
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 16206 6100 16212 6112
rect 14967 6072 16212 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 1104 6010 20700 6032
rect 1104 5958 3399 6010
rect 3451 5958 3463 6010
rect 3515 5958 3527 6010
rect 3579 5958 3591 6010
rect 3643 5958 3655 6010
rect 3707 5958 8298 6010
rect 8350 5958 8362 6010
rect 8414 5958 8426 6010
rect 8478 5958 8490 6010
rect 8542 5958 8554 6010
rect 8606 5958 13197 6010
rect 13249 5958 13261 6010
rect 13313 5958 13325 6010
rect 13377 5958 13389 6010
rect 13441 5958 13453 6010
rect 13505 5958 18096 6010
rect 18148 5958 18160 6010
rect 18212 5958 18224 6010
rect 18276 5958 18288 6010
rect 18340 5958 18352 6010
rect 18404 5958 20700 6010
rect 1104 5936 20700 5958
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 6512 5868 6561 5896
rect 6512 5856 6518 5868
rect 6549 5865 6561 5868
rect 6595 5865 6607 5899
rect 6549 5859 6607 5865
rect 9769 5899 9827 5905
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 9950 5896 9956 5908
rect 9815 5868 9956 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 13906 5896 13912 5908
rect 12207 5868 13912 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 15010 5896 15016 5908
rect 14971 5868 15016 5896
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5316 5800 6408 5828
rect 5316 5788 5322 5800
rect 3142 5760 3148 5772
rect 3103 5732 3148 5760
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 3467 5732 4261 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 6178 5760 6184 5772
rect 6139 5732 6184 5760
rect 4249 5723 4307 5729
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 6380 5769 6408 5800
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 16022 5828 16028 5840
rect 7984 5800 10456 5828
rect 15983 5800 16028 5828
rect 7984 5788 7990 5800
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 7423 5763 7481 5769
rect 7423 5729 7435 5763
rect 7469 5760 7481 5763
rect 9766 5760 9772 5772
rect 7469 5732 9772 5760
rect 7469 5729 7481 5732
rect 7423 5723 7481 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 10428 5769 10456 5800
rect 16022 5788 16028 5800
rect 16080 5788 16086 5840
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 15286 5720 15292 5772
rect 15344 5720 15350 5772
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 18598 5760 18604 5772
rect 17451 5732 18604 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 2866 5652 2872 5704
rect 2924 5692 2930 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2924 5664 3065 5692
rect 2924 5652 2930 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3053 5655 3111 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 7336 5695 7394 5701
rect 7336 5661 7348 5695
rect 7382 5692 7394 5695
rect 7382 5664 7880 5692
rect 7382 5661 7394 5664
rect 7336 5655 7394 5661
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 7852 5624 7880 5664
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 8573 5695 8631 5701
rect 7984 5664 8029 5692
rect 7984 5652 7990 5664
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8619 5664 9137 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 17126 5692 17132 5704
rect 13964 5664 15226 5692
rect 17087 5664 17132 5692
rect 13964 5652 13970 5664
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 9398 5624 9404 5636
rect 7852 5596 9404 5624
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 10689 5627 10747 5633
rect 10689 5624 10701 5627
rect 10652 5596 10701 5624
rect 10652 5584 10658 5596
rect 10689 5593 10701 5596
rect 10735 5593 10747 5627
rect 12434 5624 12440 5636
rect 11914 5596 12440 5624
rect 10689 5587 10747 5593
rect 12434 5584 12440 5596
rect 12492 5584 12498 5636
rect 19334 5624 19340 5636
rect 18630 5596 19340 5624
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5132 5528 5733 5556
rect 5132 5516 5138 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 5721 5519 5779 5525
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 17494 5556 17500 5568
rect 16439 5528 17500 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 18874 5556 18880 5568
rect 18835 5528 18880 5556
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 1104 5466 20859 5488
rect 1104 5414 5848 5466
rect 5900 5414 5912 5466
rect 5964 5414 5976 5466
rect 6028 5414 6040 5466
rect 6092 5414 6104 5466
rect 6156 5414 10747 5466
rect 10799 5414 10811 5466
rect 10863 5414 10875 5466
rect 10927 5414 10939 5466
rect 10991 5414 11003 5466
rect 11055 5414 15646 5466
rect 15698 5414 15710 5466
rect 15762 5414 15774 5466
rect 15826 5414 15838 5466
rect 15890 5414 15902 5466
rect 15954 5414 20545 5466
rect 20597 5414 20609 5466
rect 20661 5414 20673 5466
rect 20725 5414 20737 5466
rect 20789 5414 20801 5466
rect 20853 5414 20859 5466
rect 1104 5392 20859 5414
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 4706 5352 4712 5364
rect 2556 5324 4712 5352
rect 2556 5312 2562 5324
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5258 5352 5264 5364
rect 5215 5324 5264 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 6914 5352 6920 5364
rect 6875 5324 6920 5352
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 8754 5352 8760 5364
rect 7760 5324 8064 5352
rect 4724 5284 4752 5312
rect 7760 5284 7788 5324
rect 4724 5256 7788 5284
rect 4522 5216 4528 5228
rect 4483 5188 4528 5216
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 5626 5176 5632 5228
rect 5684 5225 5690 5228
rect 6748 5225 6776 5256
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 7892 5256 7941 5284
rect 7892 5244 7898 5256
rect 7929 5253 7941 5256
rect 7975 5253 7987 5287
rect 8036 5284 8064 5324
rect 8312 5324 8760 5352
rect 8312 5284 8340 5324
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9398 5352 9404 5364
rect 9359 5324 9404 5352
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 13449 5355 13507 5361
rect 12360 5324 13400 5352
rect 12360 5284 12388 5324
rect 12434 5284 12440 5296
rect 8036 5256 8418 5284
rect 12360 5256 12440 5284
rect 7929 5247 7987 5253
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 13372 5284 13400 5324
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 13906 5352 13912 5364
rect 13495 5324 13912 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14016 5324 15516 5352
rect 14016 5284 14044 5324
rect 15488 5284 15516 5324
rect 16942 5284 16948 5296
rect 13372 5256 14044 5284
rect 15410 5256 16948 5284
rect 16942 5244 16948 5256
rect 17000 5244 17006 5296
rect 17494 5284 17500 5296
rect 17455 5256 17500 5284
rect 17494 5244 17500 5256
rect 17552 5244 17558 5296
rect 19334 5284 19340 5296
rect 18722 5256 19340 5284
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 5684 5219 5722 5225
rect 5710 5185 5722 5219
rect 5684 5179 5722 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 5684 5176 5690 5179
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10045 5219 10103 5225
rect 10045 5216 10057 5219
rect 10008 5188 10057 5216
rect 10008 5176 10014 5188
rect 10045 5185 10057 5188
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 10560 5188 11713 5216
rect 10560 5176 10566 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 13872 5188 13921 5216
rect 13872 5176 13878 5188
rect 13909 5185 13921 5188
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17221 5219 17279 5225
rect 17221 5216 17233 5219
rect 17184 5188 17233 5216
rect 17184 5176 17190 5188
rect 17221 5185 17233 5188
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 7926 5148 7932 5160
rect 7699 5120 7932 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 7926 5108 7932 5120
rect 7984 5108 7990 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9861 5151 9919 5157
rect 9861 5148 9873 5151
rect 9456 5120 9873 5148
rect 9456 5108 9462 5120
rect 9861 5117 9873 5120
rect 9907 5117 9919 5151
rect 9861 5111 9919 5117
rect 10594 5108 10600 5160
rect 10652 5148 10658 5160
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 10652 5120 11989 5148
rect 10652 5108 10658 5120
rect 11977 5117 11989 5120
rect 12023 5148 12035 5151
rect 14182 5148 14188 5160
rect 12023 5120 14188 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 14182 5108 14188 5120
rect 14240 5148 14246 5160
rect 16114 5148 16120 5160
rect 14240 5120 16120 5148
rect 14240 5108 14246 5120
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 18969 5151 19027 5157
rect 18969 5117 18981 5151
rect 19015 5148 19027 5151
rect 19904 5148 19932 5179
rect 19015 5120 19932 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 5767 5083 5825 5089
rect 5767 5049 5779 5083
rect 5813 5080 5825 5083
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 5813 5052 6561 5080
rect 5813 5049 5825 5052
rect 5767 5043 5825 5049
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 6549 5043 6607 5049
rect 10226 5012 10232 5024
rect 10187 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 15657 5015 15715 5021
rect 15657 4981 15669 5015
rect 15703 5012 15715 5015
rect 15930 5012 15936 5024
rect 15703 4984 15936 5012
rect 15703 4981 15715 4984
rect 15657 4975 15715 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 20070 5012 20076 5024
rect 20031 4984 20076 5012
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 1104 4922 20700 4944
rect 1104 4870 3399 4922
rect 3451 4870 3463 4922
rect 3515 4870 3527 4922
rect 3579 4870 3591 4922
rect 3643 4870 3655 4922
rect 3707 4870 8298 4922
rect 8350 4870 8362 4922
rect 8414 4870 8426 4922
rect 8478 4870 8490 4922
rect 8542 4870 8554 4922
rect 8606 4870 13197 4922
rect 13249 4870 13261 4922
rect 13313 4870 13325 4922
rect 13377 4870 13389 4922
rect 13441 4870 13453 4922
rect 13505 4870 18096 4922
rect 18148 4870 18160 4922
rect 18212 4870 18224 4922
rect 18276 4870 18288 4922
rect 18340 4870 18352 4922
rect 18404 4870 20700 4922
rect 1104 4848 20700 4870
rect 4939 4811 4997 4817
rect 4939 4777 4951 4811
rect 4985 4808 4997 4811
rect 6178 4808 6184 4820
rect 4985 4780 6184 4808
rect 4985 4777 4997 4780
rect 4939 4771 4997 4777
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8938 4808 8944 4820
rect 8159 4780 8944 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 14921 4811 14979 4817
rect 14921 4777 14933 4811
rect 14967 4808 14979 4811
rect 16022 4808 16028 4820
rect 14967 4780 16028 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 15930 4740 15936 4752
rect 15891 4712 15936 4740
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 2832 4644 3433 4672
rect 2832 4632 2838 4644
rect 3421 4641 3433 4644
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8812 4644 9321 4672
rect 8812 4632 8818 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 9999 4675 10057 4681
rect 9999 4672 10011 4675
rect 9539 4644 10011 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 9999 4641 10011 4644
rect 10045 4641 10057 4675
rect 9999 4635 10057 4641
rect 15194 4632 15200 4684
rect 15252 4632 15258 4684
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3142 4604 3148 4616
rect 3099 4576 3148 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 4868 4607 4926 4613
rect 4868 4573 4880 4607
rect 4914 4604 4926 4607
rect 5074 4604 5080 4616
rect 4914 4576 5080 4604
rect 4914 4573 4926 4576
rect 4868 4567 4926 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 5500 4576 6377 4604
rect 5500 4564 5506 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 10102 4607 10160 4613
rect 10102 4573 10114 4607
rect 10148 4604 10160 4607
rect 10226 4604 10232 4616
rect 10148 4576 10232 4604
rect 10148 4573 10160 4576
rect 10102 4567 10160 4573
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 15378 4564 15384 4616
rect 15436 4564 15442 4616
rect 2498 4496 2504 4548
rect 2556 4496 2562 4548
rect 6638 4536 6644 4548
rect 6599 4508 6644 4536
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 7926 4536 7932 4548
rect 7839 4508 7932 4536
rect 7926 4496 7932 4508
rect 7984 4536 7990 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 7984 4508 9137 4536
rect 7984 4496 7990 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 9125 4499 9183 4505
rect 1670 4477 1676 4480
rect 1627 4471 1676 4477
rect 1627 4437 1639 4471
rect 1673 4437 1676 4471
rect 1627 4431 1676 4437
rect 1670 4428 1676 4431
rect 1728 4428 1734 4480
rect 16301 4471 16359 4477
rect 16301 4437 16313 4471
rect 16347 4468 16359 4471
rect 17678 4468 17684 4480
rect 16347 4440 17684 4468
rect 16347 4437 16359 4440
rect 16301 4431 16359 4437
rect 17678 4428 17684 4440
rect 17736 4428 17742 4480
rect 1104 4378 20859 4400
rect 1104 4326 5848 4378
rect 5900 4326 5912 4378
rect 5964 4326 5976 4378
rect 6028 4326 6040 4378
rect 6092 4326 6104 4378
rect 6156 4326 10747 4378
rect 10799 4326 10811 4378
rect 10863 4326 10875 4378
rect 10927 4326 10939 4378
rect 10991 4326 11003 4378
rect 11055 4326 15646 4378
rect 15698 4326 15710 4378
rect 15762 4326 15774 4378
rect 15826 4326 15838 4378
rect 15890 4326 15902 4378
rect 15954 4326 20545 4378
rect 20597 4326 20609 4378
rect 20661 4326 20673 4378
rect 20725 4326 20737 4378
rect 20789 4326 20801 4378
rect 20853 4326 20859 4378
rect 1104 4304 20859 4326
rect 6638 4273 6644 4276
rect 6595 4267 6644 4273
rect 6595 4233 6607 4267
rect 6641 4233 6644 4267
rect 6595 4227 6644 4233
rect 6638 4224 6644 4227
rect 6696 4224 6702 4276
rect 2498 4156 2504 4208
rect 2556 4156 2562 4208
rect 8754 4156 8760 4208
rect 8812 4156 8818 4208
rect 19334 4196 19340 4208
rect 19274 4168 19340 4196
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 3200 4100 3249 4128
rect 3200 4088 3206 4100
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 6454 4128 6460 4140
rect 3651 4100 6460 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6698 4131 6756 4137
rect 6698 4097 6710 4131
rect 6744 4128 6756 4131
rect 8021 4131 8079 4137
rect 6744 4097 6776 4128
rect 6698 4091 6776 4097
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8067 4100 8524 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 6748 4060 6776 4091
rect 7374 4060 7380 4072
rect 6748 4032 7380 4060
rect 7374 4020 7380 4032
rect 7432 4060 7438 4072
rect 8202 4060 8208 4072
rect 7432 4032 8208 4060
rect 7432 4020 7438 4032
rect 8202 4020 8208 4032
rect 8260 4060 8266 4072
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8260 4032 8401 4060
rect 8260 4020 8266 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8496 4060 8524 4100
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17184 4100 17785 4128
rect 17184 4088 17190 4100
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 10410 4060 10416 4072
rect 8496 4032 10416 4060
rect 8389 4023 8447 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17880 4032 18061 4060
rect 17678 3952 17684 4004
rect 17736 3992 17742 4004
rect 17880 3992 17908 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 17736 3964 17908 3992
rect 17736 3952 17742 3964
rect 1811 3927 1869 3933
rect 1811 3893 1823 3927
rect 1857 3924 1869 3927
rect 2314 3924 2320 3936
rect 1857 3896 2320 3924
rect 1857 3893 1869 3896
rect 1811 3887 1869 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 9674 3924 9680 3936
rect 3016 3896 9680 3924
rect 3016 3884 3022 3896
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 9815 3927 9873 3933
rect 9815 3893 9827 3927
rect 9861 3924 9873 3927
rect 9950 3924 9956 3936
rect 9861 3896 9956 3924
rect 9861 3893 9873 3896
rect 9815 3887 9873 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 19521 3927 19579 3933
rect 19521 3893 19533 3927
rect 19567 3924 19579 3927
rect 19886 3924 19892 3936
rect 19567 3896 19892 3924
rect 19567 3893 19579 3896
rect 19521 3887 19579 3893
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 1104 3834 20700 3856
rect 1104 3782 3399 3834
rect 3451 3782 3463 3834
rect 3515 3782 3527 3834
rect 3579 3782 3591 3834
rect 3643 3782 3655 3834
rect 3707 3782 8298 3834
rect 8350 3782 8362 3834
rect 8414 3782 8426 3834
rect 8478 3782 8490 3834
rect 8542 3782 8554 3834
rect 8606 3782 13197 3834
rect 13249 3782 13261 3834
rect 13313 3782 13325 3834
rect 13377 3782 13389 3834
rect 13441 3782 13453 3834
rect 13505 3782 18096 3834
rect 18148 3782 18160 3834
rect 18212 3782 18224 3834
rect 18276 3782 18288 3834
rect 18340 3782 18352 3834
rect 18404 3782 20700 3834
rect 1104 3760 20700 3782
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 2409 3655 2467 3661
rect 2409 3652 2421 3655
rect 624 3624 2421 3652
rect 624 3612 630 3624
rect 2409 3621 2421 3624
rect 2455 3621 2467 3655
rect 2409 3615 2467 3621
rect 10594 3612 10600 3664
rect 10652 3612 10658 3664
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 4304 3556 5089 3584
rect 4304 3544 4310 3556
rect 5077 3553 5089 3556
rect 5123 3584 5135 3587
rect 5442 3584 5448 3596
rect 5123 3556 5448 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 10612 3584 10640 3612
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10612 3556 10977 3584
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 11514 3584 11520 3596
rect 10965 3547 11023 3553
rect 11072 3556 11520 3584
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 3234 3516 3240 3528
rect 2639 3488 3240 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 11072 3516 11100 3556
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3584 15899 3587
rect 16022 3584 16028 3596
rect 15887 3556 16028 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 19886 3516 19892 3528
rect 10643 3488 11100 3516
rect 19847 3488 19892 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 5350 3448 5356 3460
rect 5311 3420 5356 3448
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 6914 3448 6920 3460
rect 6578 3420 6920 3448
rect 6914 3408 6920 3420
rect 6972 3408 6978 3460
rect 11330 3408 11336 3460
rect 11388 3408 11394 3460
rect 16850 3408 16856 3460
rect 16908 3408 16914 3460
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 4430 3380 4436 3392
rect 4391 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 6825 3383 6883 3389
rect 6825 3349 6837 3383
rect 6871 3380 6883 3383
rect 7098 3380 7104 3392
rect 6871 3352 7104 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 12391 3383 12449 3389
rect 12391 3349 12403 3383
rect 12437 3380 12449 3383
rect 12526 3380 12532 3392
rect 12437 3352 12532 3380
rect 12437 3349 12449 3352
rect 12391 3343 12449 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 17267 3383 17325 3389
rect 17267 3349 17279 3383
rect 17313 3380 17325 3383
rect 17402 3380 17408 3392
rect 17313 3352 17408 3380
rect 17313 3349 17325 3352
rect 17267 3343 17325 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 20070 3380 20076 3392
rect 20031 3352 20076 3380
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 1104 3290 20859 3312
rect 1104 3238 5848 3290
rect 5900 3238 5912 3290
rect 5964 3238 5976 3290
rect 6028 3238 6040 3290
rect 6092 3238 6104 3290
rect 6156 3238 10747 3290
rect 10799 3238 10811 3290
rect 10863 3238 10875 3290
rect 10927 3238 10939 3290
rect 10991 3238 11003 3290
rect 11055 3238 15646 3290
rect 15698 3238 15710 3290
rect 15762 3238 15774 3290
rect 15826 3238 15838 3290
rect 15890 3238 15902 3290
rect 15954 3238 20545 3290
rect 20597 3238 20609 3290
rect 20661 3238 20673 3290
rect 20725 3238 20737 3290
rect 20789 3238 20801 3290
rect 20853 3238 20859 3290
rect 1104 3216 20859 3238
rect 2498 3136 2504 3188
rect 2556 3176 2562 3188
rect 2556 3148 3740 3176
rect 2556 3136 2562 3148
rect 3712 3108 3740 3148
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4847 3179 4905 3185
rect 4847 3176 4859 3179
rect 4672 3148 4859 3176
rect 4672 3136 4678 3148
rect 4847 3145 4859 3148
rect 4893 3145 4905 3179
rect 4847 3139 4905 3145
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 16908 3148 17540 3176
rect 16908 3136 16914 3148
rect 3712 3080 3818 3108
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 6825 3111 6883 3117
rect 6825 3108 6837 3111
rect 5408 3080 6837 3108
rect 5408 3068 5414 3080
rect 6825 3077 6837 3080
rect 6871 3077 6883 3111
rect 11330 3108 11336 3120
rect 10718 3080 11336 3108
rect 6825 3071 6883 3077
rect 11330 3068 11336 3080
rect 11388 3108 11394 3120
rect 12434 3108 12440 3120
rect 11388 3080 12440 3108
rect 11388 3068 11394 3080
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 17512 3108 17540 3148
rect 17512 3080 17618 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 1670 3040 1676 3052
rect 1627 3012 1676 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 3016 3012 3065 3040
rect 3016 3000 3022 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3200 3012 3433 3040
rect 3200 3000 3206 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 5994 3040 6000 3052
rect 5955 3012 6000 3040
rect 3421 3003 3479 3009
rect 3436 2972 3464 3003
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 7926 3000 7932 3052
rect 7984 3000 7990 3052
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9766 3040 9772 3052
rect 9355 3012 9772 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16816 3012 16865 3040
rect 16816 3000 16822 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 18932 3012 19165 3040
rect 18932 3000 18938 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 19794 3000 19800 3052
rect 19852 3040 19858 3052
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19852 3012 19901 3040
rect 19852 3000 19858 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 3786 2972 3792 2984
rect 3436 2944 3792 2972
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 4304 2944 6561 2972
rect 4304 2932 4310 2944
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 8260 2944 9689 2972
rect 8260 2932 8266 2944
rect 9677 2941 9689 2944
rect 9723 2941 9735 2975
rect 9677 2935 9735 2941
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 16080 2944 17233 2972
rect 16080 2932 16086 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 18647 2975 18705 2981
rect 18647 2941 18659 2975
rect 18693 2972 18705 2975
rect 19426 2972 19432 2984
rect 18693 2944 19432 2972
rect 18693 2941 18705 2944
rect 18647 2935 18705 2941
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 21174 2904 21180 2916
rect 19300 2876 21180 2904
rect 19300 2864 19306 2876
rect 21174 2864 21180 2876
rect 21232 2864 21238 2916
rect 1765 2839 1823 2845
rect 1765 2805 1777 2839
rect 1811 2836 1823 2839
rect 1854 2836 1860 2848
rect 1811 2808 1860 2836
rect 1811 2805 1823 2808
rect 1765 2799 1823 2805
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 2501 2839 2559 2845
rect 2501 2805 2513 2839
rect 2547 2836 2559 2839
rect 3050 2836 3056 2848
rect 2547 2808 3056 2836
rect 2547 2805 2559 2808
rect 2501 2799 2559 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 5813 2839 5871 2845
rect 5813 2836 5825 2839
rect 5776 2808 5825 2836
rect 5776 2796 5782 2808
rect 5813 2805 5825 2808
rect 5859 2805 5871 2839
rect 5813 2799 5871 2805
rect 8297 2839 8355 2845
rect 8297 2805 8309 2839
rect 8343 2836 8355 2839
rect 8662 2836 8668 2848
rect 8343 2808 8668 2836
rect 8343 2805 8355 2808
rect 8297 2799 8355 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 11146 2845 11152 2848
rect 11103 2839 11152 2845
rect 11103 2805 11115 2839
rect 11149 2805 11152 2839
rect 11103 2799 11152 2805
rect 11146 2796 11152 2799
rect 11204 2796 11210 2848
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19337 2839 19395 2845
rect 19337 2836 19349 2839
rect 19208 2808 19349 2836
rect 19208 2796 19214 2808
rect 19337 2805 19349 2808
rect 19383 2805 19395 2839
rect 19337 2799 19395 2805
rect 19886 2796 19892 2848
rect 19944 2836 19950 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 19944 2808 20085 2836
rect 19944 2796 19950 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 1104 2746 20700 2768
rect 1104 2694 3399 2746
rect 3451 2694 3463 2746
rect 3515 2694 3527 2746
rect 3579 2694 3591 2746
rect 3643 2694 3655 2746
rect 3707 2694 8298 2746
rect 8350 2694 8362 2746
rect 8414 2694 8426 2746
rect 8478 2694 8490 2746
rect 8542 2694 8554 2746
rect 8606 2694 13197 2746
rect 13249 2694 13261 2746
rect 13313 2694 13325 2746
rect 13377 2694 13389 2746
rect 13441 2694 13453 2746
rect 13505 2694 18096 2746
rect 18148 2694 18160 2746
rect 18212 2694 18224 2746
rect 18276 2694 18288 2746
rect 18340 2694 18352 2746
rect 18404 2694 20700 2746
rect 1104 2672 20700 2694
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 3292 2604 3341 2632
rect 3292 2592 3298 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 3329 2595 3387 2601
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 4328 2635 4386 2641
rect 4328 2632 4340 2635
rect 3844 2604 4340 2632
rect 3844 2592 3850 2604
rect 4328 2601 4340 2604
rect 4374 2632 4386 2635
rect 5350 2632 5356 2644
rect 4374 2604 5356 2632
rect 4374 2601 4386 2604
rect 4328 2595 4386 2601
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 5994 2632 6000 2644
rect 5859 2604 6000 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 18693 2635 18751 2641
rect 18693 2601 18705 2635
rect 18739 2632 18751 2635
rect 19242 2632 19248 2644
rect 18739 2604 19248 2632
rect 18739 2601 18751 2604
rect 18693 2595 18751 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 9490 2496 9496 2508
rect 1627 2468 9496 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 19702 2496 19708 2508
rect 18892 2468 19708 2496
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 7098 2428 7104 2440
rect 7059 2400 7104 2428
rect 4065 2391 4123 2397
rect 1857 2363 1915 2369
rect 1857 2329 1869 2363
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 1872 2292 1900 2323
rect 2498 2320 2504 2372
rect 2556 2320 2562 2372
rect 4080 2360 4108 2391
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8662 2428 8668 2440
rect 8343 2400 8668 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 11146 2428 11152 2440
rect 11107 2400 11152 2428
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 12526 2428 12532 2440
rect 12487 2400 12532 2428
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 14274 2428 14280 2440
rect 14235 2400 14280 2428
rect 14274 2388 14280 2400
rect 14332 2388 14338 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15378 2428 15384 2440
rect 15335 2400 15384 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16724 2400 16865 2428
rect 16724 2388 16730 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 18892 2437 18920 2468
rect 19702 2456 19708 2468
rect 19760 2456 19766 2508
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17460 2400 17601 2428
rect 17460 2388 17466 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 18877 2391 18935 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 4246 2360 4252 2372
rect 4080 2332 4252 2360
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 4798 2320 4804 2372
rect 4856 2320 4862 2372
rect 3786 2292 3792 2304
rect 1872 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7064 2264 7297 2292
rect 7064 2252 7070 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8352 2264 8493 2292
rect 8352 2252 8358 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9640 2264 9781 2292
rect 9640 2252 9646 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 10965 2295 11023 2301
rect 10965 2292 10977 2295
rect 10652 2264 10977 2292
rect 10652 2252 10658 2264
rect 10965 2261 10977 2264
rect 11011 2261 11023 2295
rect 10965 2255 11023 2261
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12216 2264 12357 2292
rect 12216 2252 12222 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 13504 2264 14473 2292
rect 13504 2252 13510 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14792 2264 15117 2292
rect 14792 2252 14798 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16080 2264 17049 2292
rect 16080 2252 16086 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 17773 2295 17831 2301
rect 17773 2292 17785 2295
rect 17368 2264 17785 2292
rect 17368 2252 17374 2264
rect 17773 2261 17785 2264
rect 17819 2261 17831 2295
rect 17773 2255 17831 2261
rect 18874 2252 18880 2304
rect 18932 2292 18938 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 18932 2264 19625 2292
rect 18932 2252 18938 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 1104 2202 20859 2224
rect 1104 2150 5848 2202
rect 5900 2150 5912 2202
rect 5964 2150 5976 2202
rect 6028 2150 6040 2202
rect 6092 2150 6104 2202
rect 6156 2150 10747 2202
rect 10799 2150 10811 2202
rect 10863 2150 10875 2202
rect 10927 2150 10939 2202
rect 10991 2150 11003 2202
rect 11055 2150 15646 2202
rect 15698 2150 15710 2202
rect 15762 2150 15774 2202
rect 15826 2150 15838 2202
rect 15890 2150 15902 2202
rect 15954 2150 20545 2202
rect 20597 2150 20609 2202
rect 20661 2150 20673 2202
rect 20725 2150 20737 2202
rect 20789 2150 20801 2202
rect 20853 2150 20859 2202
rect 1104 2128 20859 2150
<< via1 >>
rect 5848 21734 5900 21786
rect 5912 21734 5964 21786
rect 5976 21734 6028 21786
rect 6040 21734 6092 21786
rect 6104 21734 6156 21786
rect 10747 21734 10799 21786
rect 10811 21734 10863 21786
rect 10875 21734 10927 21786
rect 10939 21734 10991 21786
rect 11003 21734 11055 21786
rect 15646 21734 15698 21786
rect 15710 21734 15762 21786
rect 15774 21734 15826 21786
rect 15838 21734 15890 21786
rect 15902 21734 15954 21786
rect 20545 21734 20597 21786
rect 20609 21734 20661 21786
rect 20673 21734 20725 21786
rect 20737 21734 20789 21786
rect 20801 21734 20853 21786
rect 1860 21632 1912 21684
rect 3148 21632 3200 21684
rect 4620 21675 4672 21684
rect 4620 21641 4629 21675
rect 4629 21641 4663 21675
rect 4663 21641 4672 21675
rect 4620 21632 4672 21641
rect 5724 21632 5776 21684
rect 7288 21675 7340 21684
rect 7288 21641 7297 21675
rect 7297 21641 7331 21675
rect 7331 21641 7340 21675
rect 7288 21632 7340 21641
rect 8300 21632 8352 21684
rect 9680 21632 9732 21684
rect 10600 21632 10652 21684
rect 12348 21675 12400 21684
rect 12348 21641 12357 21675
rect 12357 21641 12391 21675
rect 12391 21641 12400 21675
rect 12348 21632 12400 21641
rect 13820 21632 13872 21684
rect 14740 21632 14792 21684
rect 16028 21632 16080 21684
rect 17316 21632 17368 21684
rect 18604 21632 18656 21684
rect 3240 21496 3292 21548
rect 4068 21496 4120 21548
rect 4896 21496 4948 21548
rect 5632 21496 5684 21548
rect 7472 21496 7524 21548
rect 8944 21496 8996 21548
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 12532 21539 12584 21548
rect 12532 21505 12541 21539
rect 12541 21505 12575 21539
rect 12575 21505 12584 21539
rect 12532 21496 12584 21505
rect 14188 21496 14240 21548
rect 14372 21496 14424 21548
rect 16580 21496 16632 21548
rect 17592 21539 17644 21548
rect 17592 21505 17601 21539
rect 17601 21505 17635 21539
rect 17635 21505 17644 21539
rect 17592 21496 17644 21505
rect 18880 21539 18932 21548
rect 18880 21505 18889 21539
rect 18889 21505 18923 21539
rect 18923 21505 18932 21539
rect 18880 21496 18932 21505
rect 19064 21496 19116 21548
rect 16672 21428 16724 21480
rect 21180 21360 21232 21412
rect 15752 21292 15804 21344
rect 3399 21190 3451 21242
rect 3463 21190 3515 21242
rect 3527 21190 3579 21242
rect 3591 21190 3643 21242
rect 3655 21190 3707 21242
rect 8298 21190 8350 21242
rect 8362 21190 8414 21242
rect 8426 21190 8478 21242
rect 8490 21190 8542 21242
rect 8554 21190 8606 21242
rect 13197 21190 13249 21242
rect 13261 21190 13313 21242
rect 13325 21190 13377 21242
rect 13389 21190 13441 21242
rect 13453 21190 13505 21242
rect 18096 21190 18148 21242
rect 18160 21190 18212 21242
rect 18224 21190 18276 21242
rect 18288 21190 18340 21242
rect 18352 21190 18404 21242
rect 572 21088 624 21140
rect 14280 21088 14332 21140
rect 17592 21088 17644 21140
rect 19892 21088 19944 21140
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 2688 20927 2740 20936
rect 2688 20893 2697 20927
rect 2697 20893 2731 20927
rect 2731 20893 2740 20927
rect 2688 20884 2740 20893
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 15752 20995 15804 21004
rect 6552 20884 6604 20893
rect 9496 20884 9548 20936
rect 10140 20927 10192 20936
rect 10140 20893 10149 20927
rect 10149 20893 10183 20927
rect 10183 20893 10192 20927
rect 10140 20884 10192 20893
rect 13452 20927 13504 20936
rect 13452 20893 13461 20927
rect 13461 20893 13495 20927
rect 13495 20893 13504 20927
rect 13452 20884 13504 20893
rect 15292 20884 15344 20936
rect 15752 20961 15761 20995
rect 15761 20961 15795 20995
rect 15795 20961 15804 20995
rect 15752 20952 15804 20961
rect 19248 20952 19300 21004
rect 16672 20884 16724 20936
rect 18420 20927 18472 20936
rect 18420 20893 18454 20927
rect 18454 20893 18472 20927
rect 19892 20927 19944 20936
rect 18420 20884 18472 20893
rect 19892 20893 19901 20927
rect 19901 20893 19935 20927
rect 19935 20893 19944 20927
rect 19892 20884 19944 20893
rect 2780 20816 2832 20868
rect 3884 20816 3936 20868
rect 6920 20816 6972 20868
rect 10416 20859 10468 20868
rect 10416 20825 10425 20859
rect 10425 20825 10459 20859
rect 10459 20825 10468 20859
rect 10416 20816 10468 20825
rect 11428 20816 11480 20868
rect 17592 20816 17644 20868
rect 5540 20748 5592 20800
rect 8300 20748 8352 20800
rect 11336 20748 11388 20800
rect 17224 20748 17276 20800
rect 17868 20748 17920 20800
rect 5848 20646 5900 20698
rect 5912 20646 5964 20698
rect 5976 20646 6028 20698
rect 6040 20646 6092 20698
rect 6104 20646 6156 20698
rect 10747 20646 10799 20698
rect 10811 20646 10863 20698
rect 10875 20646 10927 20698
rect 10939 20646 10991 20698
rect 11003 20646 11055 20698
rect 15646 20646 15698 20698
rect 15710 20646 15762 20698
rect 15774 20646 15826 20698
rect 15838 20646 15890 20698
rect 15902 20646 15954 20698
rect 20545 20646 20597 20698
rect 20609 20646 20661 20698
rect 20673 20646 20725 20698
rect 20737 20646 20789 20698
rect 20801 20646 20853 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 9680 20544 9732 20596
rect 2780 20476 2832 20528
rect 4252 20476 4304 20528
rect 9864 20476 9916 20528
rect 13452 20544 13504 20596
rect 19064 20544 19116 20596
rect 19248 20587 19300 20596
rect 19248 20553 19257 20587
rect 19257 20553 19291 20587
rect 19291 20553 19300 20587
rect 19248 20544 19300 20553
rect 2596 20451 2648 20460
rect 2596 20417 2605 20451
rect 2605 20417 2639 20451
rect 2639 20417 2648 20451
rect 2596 20408 2648 20417
rect 7288 20408 7340 20460
rect 8024 20408 8076 20460
rect 8300 20451 8352 20460
rect 8300 20417 8309 20451
rect 8309 20417 8343 20451
rect 8343 20417 8352 20451
rect 8300 20408 8352 20417
rect 10140 20408 10192 20460
rect 11060 20408 11112 20460
rect 17592 20476 17644 20528
rect 5724 20340 5776 20392
rect 10324 20340 10376 20392
rect 12808 20340 12860 20392
rect 2780 20247 2832 20256
rect 2780 20213 2789 20247
rect 2789 20213 2823 20247
rect 2823 20213 2832 20247
rect 2780 20204 2832 20213
rect 4252 20204 4304 20256
rect 7012 20204 7064 20256
rect 12440 20204 12492 20256
rect 15384 20408 15436 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 19524 20408 19576 20460
rect 13452 20340 13504 20392
rect 16028 20340 16080 20392
rect 16764 20340 16816 20392
rect 15476 20204 15528 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 3399 20102 3451 20154
rect 3463 20102 3515 20154
rect 3527 20102 3579 20154
rect 3591 20102 3643 20154
rect 3655 20102 3707 20154
rect 8298 20102 8350 20154
rect 8362 20102 8414 20154
rect 8426 20102 8478 20154
rect 8490 20102 8542 20154
rect 8554 20102 8606 20154
rect 13197 20102 13249 20154
rect 13261 20102 13313 20154
rect 13325 20102 13377 20154
rect 13389 20102 13441 20154
rect 13453 20102 13505 20154
rect 18096 20102 18148 20154
rect 18160 20102 18212 20154
rect 18224 20102 18276 20154
rect 18288 20102 18340 20154
rect 18352 20102 18404 20154
rect 2688 20000 2740 20052
rect 7288 20000 7340 20052
rect 12808 20043 12860 20052
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 5540 19864 5592 19916
rect 9220 19864 9272 19916
rect 11060 19907 11112 19916
rect 11060 19873 11069 19907
rect 11069 19873 11103 19907
rect 11103 19873 11112 19907
rect 11060 19864 11112 19873
rect 11336 19907 11388 19916
rect 11336 19873 11345 19907
rect 11345 19873 11379 19907
rect 11379 19873 11388 19907
rect 11336 19864 11388 19873
rect 15752 19907 15804 19916
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 16028 19907 16080 19916
rect 16028 19873 16037 19907
rect 16037 19873 16071 19907
rect 16071 19873 16080 19907
rect 16028 19864 16080 19873
rect 17868 19864 17920 19916
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 2780 19796 2832 19805
rect 5724 19796 5776 19848
rect 12440 19796 12492 19848
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 17132 19839 17184 19848
rect 17132 19805 17141 19839
rect 17141 19805 17175 19839
rect 17175 19805 17184 19839
rect 17132 19796 17184 19805
rect 18880 19796 18932 19848
rect 6552 19728 6604 19780
rect 7012 19728 7064 19780
rect 15476 19728 15528 19780
rect 17040 19728 17092 19780
rect 18972 19728 19024 19780
rect 8024 19660 8076 19712
rect 11244 19660 11296 19712
rect 18696 19660 18748 19712
rect 5848 19558 5900 19610
rect 5912 19558 5964 19610
rect 5976 19558 6028 19610
rect 6040 19558 6092 19610
rect 6104 19558 6156 19610
rect 10747 19558 10799 19610
rect 10811 19558 10863 19610
rect 10875 19558 10927 19610
rect 10939 19558 10991 19610
rect 11003 19558 11055 19610
rect 15646 19558 15698 19610
rect 15710 19558 15762 19610
rect 15774 19558 15826 19610
rect 15838 19558 15890 19610
rect 15902 19558 15954 19610
rect 20545 19558 20597 19610
rect 20609 19558 20661 19610
rect 20673 19558 20725 19610
rect 20737 19558 20789 19610
rect 20801 19558 20853 19610
rect 2596 19431 2648 19440
rect 2596 19397 2605 19431
rect 2605 19397 2639 19431
rect 2639 19397 2648 19431
rect 2596 19388 2648 19397
rect 4252 19388 4304 19440
rect 8024 19388 8076 19440
rect 10416 19456 10468 19508
rect 19432 19456 19484 19508
rect 11244 19388 11296 19440
rect 18972 19388 19024 19440
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 16212 19320 16264 19372
rect 17868 19320 17920 19372
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 17132 19252 17184 19304
rect 17960 19252 18012 19304
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 4252 19116 4304 19168
rect 8668 19116 8720 19168
rect 17224 19116 17276 19168
rect 19708 19116 19760 19168
rect 3399 19014 3451 19066
rect 3463 19014 3515 19066
rect 3527 19014 3579 19066
rect 3591 19014 3643 19066
rect 3655 19014 3707 19066
rect 8298 19014 8350 19066
rect 8362 19014 8414 19066
rect 8426 19014 8478 19066
rect 8490 19014 8542 19066
rect 8554 19014 8606 19066
rect 13197 19014 13249 19066
rect 13261 19014 13313 19066
rect 13325 19014 13377 19066
rect 13389 19014 13441 19066
rect 13453 19014 13505 19066
rect 18096 19014 18148 19066
rect 18160 19014 18212 19066
rect 18224 19014 18276 19066
rect 18288 19014 18340 19066
rect 18352 19014 18404 19066
rect 8668 18912 8720 18964
rect 12532 18912 12584 18964
rect 17868 18955 17920 18964
rect 17868 18921 17877 18955
rect 17877 18921 17911 18955
rect 17911 18921 17920 18955
rect 17868 18912 17920 18921
rect 17040 18844 17092 18896
rect 19800 18844 19852 18896
rect 2320 18776 2372 18828
rect 4252 18819 4304 18828
rect 4252 18785 4261 18819
rect 4261 18785 4295 18819
rect 4295 18785 4304 18819
rect 4252 18776 4304 18785
rect 12440 18776 12492 18828
rect 16212 18776 16264 18828
rect 6552 18708 6604 18760
rect 4344 18640 4396 18692
rect 7104 18683 7156 18692
rect 7104 18649 7113 18683
rect 7113 18649 7147 18683
rect 7147 18649 7156 18683
rect 7104 18640 7156 18649
rect 5080 18572 5132 18624
rect 5632 18572 5684 18624
rect 7012 18572 7064 18624
rect 7564 18640 7616 18692
rect 15384 18708 15436 18760
rect 17040 18751 17092 18760
rect 17040 18717 17049 18751
rect 17049 18717 17083 18751
rect 17083 18717 17092 18751
rect 17040 18708 17092 18717
rect 18512 18751 18564 18760
rect 18512 18717 18520 18751
rect 18520 18717 18564 18751
rect 18512 18708 18564 18717
rect 20260 18708 20312 18760
rect 12072 18640 12124 18692
rect 16028 18640 16080 18692
rect 11704 18572 11756 18624
rect 18144 18572 18196 18624
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 1120 18460 1470 18540
rect 5848 18470 5900 18522
rect 5912 18470 5964 18522
rect 5976 18470 6028 18522
rect 6040 18470 6092 18522
rect 6104 18470 6156 18522
rect 10747 18470 10799 18522
rect 10811 18470 10863 18522
rect 10875 18470 10927 18522
rect 10939 18470 10991 18522
rect 11003 18470 11055 18522
rect 15646 18470 15698 18522
rect 15710 18470 15762 18522
rect 15774 18470 15826 18522
rect 15838 18470 15890 18522
rect 15902 18470 15954 18522
rect 20545 18470 20597 18522
rect 20609 18470 20661 18522
rect 20673 18470 20725 18522
rect 20737 18470 20789 18522
rect 20801 18470 20853 18522
rect 7012 18368 7064 18420
rect 7104 18368 7156 18420
rect 11152 18368 11204 18420
rect 12440 18368 12492 18420
rect 5632 18343 5684 18352
rect 5632 18309 5641 18343
rect 5641 18309 5675 18343
rect 5675 18309 5684 18343
rect 5632 18300 5684 18309
rect 7564 18300 7616 18352
rect 12072 18300 12124 18352
rect 2320 18232 2372 18284
rect 4528 18232 4580 18284
rect 5080 18164 5132 18216
rect 6552 18207 6604 18216
rect 6552 18173 6561 18207
rect 6561 18173 6595 18207
rect 6595 18173 6604 18207
rect 6552 18164 6604 18173
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 10232 18164 10284 18216
rect 12440 18232 12492 18284
rect 15384 18368 15436 18420
rect 16212 18411 16264 18420
rect 16212 18377 16221 18411
rect 16221 18377 16255 18411
rect 16255 18377 16264 18411
rect 16212 18368 16264 18377
rect 16028 18300 16080 18352
rect 18880 18368 18932 18420
rect 19892 18368 19944 18420
rect 18144 18343 18196 18352
rect 18144 18309 18153 18343
rect 18153 18309 18187 18343
rect 18187 18309 18196 18343
rect 18144 18300 18196 18309
rect 18788 18300 18840 18352
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 14280 18164 14332 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 17868 18207 17920 18216
rect 17868 18173 17877 18207
rect 17877 18173 17911 18207
rect 17911 18173 17920 18207
rect 17868 18164 17920 18173
rect 1952 18028 2004 18080
rect 4160 18071 4212 18080
rect 4160 18037 4169 18071
rect 4169 18037 4203 18071
rect 4203 18037 4212 18071
rect 4160 18028 4212 18037
rect 12440 18028 12492 18080
rect 16764 18028 16816 18080
rect 3399 17926 3451 17978
rect 3463 17926 3515 17978
rect 3527 17926 3579 17978
rect 3591 17926 3643 17978
rect 3655 17926 3707 17978
rect 8298 17926 8350 17978
rect 8362 17926 8414 17978
rect 8426 17926 8478 17978
rect 8490 17926 8542 17978
rect 8554 17926 8606 17978
rect 13197 17926 13249 17978
rect 13261 17926 13313 17978
rect 13325 17926 13377 17978
rect 13389 17926 13441 17978
rect 13453 17926 13505 17978
rect 18096 17926 18148 17978
rect 18160 17926 18212 17978
rect 18224 17926 18276 17978
rect 18288 17926 18340 17978
rect 18352 17926 18404 17978
rect 6828 17867 6880 17876
rect 6828 17833 6837 17867
rect 6837 17833 6871 17867
rect 6871 17833 6880 17867
rect 6828 17824 6880 17833
rect 9680 17824 9732 17876
rect 11244 17824 11296 17876
rect 14740 17824 14792 17876
rect 19524 17824 19576 17876
rect 4160 17688 4212 17740
rect 12440 17688 12492 17740
rect 14096 17688 14148 17740
rect 14280 17688 14332 17740
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 17776 17731 17828 17740
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 1952 17663 2004 17672
rect 1952 17629 1961 17663
rect 1961 17629 1995 17663
rect 1995 17629 2004 17663
rect 1952 17620 2004 17629
rect 2688 17620 2740 17672
rect 5080 17663 5132 17672
rect 2504 17484 2556 17536
rect 3056 17484 3108 17536
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 9496 17663 9548 17672
rect 4528 17552 4580 17604
rect 9496 17629 9540 17663
rect 9540 17629 9548 17663
rect 9496 17620 9548 17629
rect 13728 17663 13780 17672
rect 9680 17552 9732 17604
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 17684 17620 17736 17672
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 7932 17484 7984 17536
rect 17776 17552 17828 17604
rect 19800 17552 19852 17604
rect 20076 17595 20128 17604
rect 20076 17561 20085 17595
rect 20085 17561 20119 17595
rect 20119 17561 20128 17595
rect 20076 17552 20128 17561
rect 17868 17484 17920 17536
rect 18604 17484 18656 17536
rect 5848 17382 5900 17434
rect 5912 17382 5964 17434
rect 5976 17382 6028 17434
rect 6040 17382 6092 17434
rect 6104 17382 6156 17434
rect 10747 17382 10799 17434
rect 10811 17382 10863 17434
rect 10875 17382 10927 17434
rect 10939 17382 10991 17434
rect 11003 17382 11055 17434
rect 15646 17382 15698 17434
rect 15710 17382 15762 17434
rect 15774 17382 15826 17434
rect 15838 17382 15890 17434
rect 15902 17382 15954 17434
rect 20545 17382 20597 17434
rect 20609 17382 20661 17434
rect 20673 17382 20725 17434
rect 20737 17382 20789 17434
rect 20801 17382 20853 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 15384 17280 15436 17332
rect 16488 17280 16540 17332
rect 17592 17280 17644 17332
rect 2596 17212 2648 17264
rect 3056 17255 3108 17264
rect 3056 17221 3065 17255
rect 3065 17221 3099 17255
rect 3099 17221 3108 17255
rect 3056 17212 3108 17221
rect 3148 17212 3200 17264
rect 18604 17212 18656 17264
rect 3884 17187 3936 17196
rect 3884 17153 3902 17187
rect 3902 17153 3936 17187
rect 3884 17144 3936 17153
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 9496 17187 9548 17196
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 14648 17187 14700 17196
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 17868 17187 17920 17196
rect 17868 17153 17877 17187
rect 17877 17153 17911 17187
rect 17911 17153 17920 17187
rect 17868 17144 17920 17153
rect 15476 17076 15528 17128
rect 17500 17076 17552 17128
rect 18512 17076 18564 17128
rect 16028 17008 16080 17060
rect 3976 16940 4028 16992
rect 6828 16940 6880 16992
rect 7748 16983 7800 16992
rect 7748 16949 7757 16983
rect 7757 16949 7791 16983
rect 7791 16949 7800 16983
rect 7748 16940 7800 16949
rect 19892 16940 19944 16992
rect 3399 16838 3451 16890
rect 3463 16838 3515 16890
rect 3527 16838 3579 16890
rect 3591 16838 3643 16890
rect 3655 16838 3707 16890
rect 8298 16838 8350 16890
rect 8362 16838 8414 16890
rect 8426 16838 8478 16890
rect 8490 16838 8542 16890
rect 8554 16838 8606 16890
rect 13197 16838 13249 16890
rect 13261 16838 13313 16890
rect 13325 16838 13377 16890
rect 13389 16838 13441 16890
rect 13453 16838 13505 16890
rect 18096 16838 18148 16890
rect 18160 16838 18212 16890
rect 18224 16838 18276 16890
rect 18288 16838 18340 16890
rect 18352 16838 18404 16890
rect 8668 16736 8720 16788
rect 9496 16736 9548 16788
rect 12532 16736 12584 16788
rect 16028 16779 16080 16788
rect 2044 16600 2096 16652
rect 2504 16643 2556 16652
rect 2504 16609 2513 16643
rect 2513 16609 2547 16643
rect 2547 16609 2556 16643
rect 2504 16600 2556 16609
rect 3976 16643 4028 16652
rect 3976 16609 3985 16643
rect 3985 16609 4019 16643
rect 4019 16609 4028 16643
rect 3976 16600 4028 16609
rect 3884 16532 3936 16584
rect 4528 16600 4580 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7748 16600 7800 16652
rect 10416 16600 10468 16652
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 12440 16600 12492 16652
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16488 16643 16540 16652
rect 16488 16609 16497 16643
rect 16497 16609 16531 16643
rect 16531 16609 16540 16643
rect 16488 16600 16540 16609
rect 17500 16600 17552 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 20168 16575 20220 16584
rect 20168 16541 20177 16575
rect 20177 16541 20211 16575
rect 20211 16541 20220 16575
rect 20168 16532 20220 16541
rect 8116 16464 8168 16516
rect 9772 16464 9824 16516
rect 13728 16464 13780 16516
rect 15936 16464 15988 16516
rect 16120 16464 16172 16516
rect 17776 16464 17828 16516
rect 5632 16396 5684 16448
rect 11612 16396 11664 16448
rect 18512 16396 18564 16448
rect 19984 16439 20036 16448
rect 19984 16405 19993 16439
rect 19993 16405 20027 16439
rect 20027 16405 20036 16439
rect 19984 16396 20036 16405
rect 5848 16294 5900 16346
rect 5912 16294 5964 16346
rect 5976 16294 6028 16346
rect 6040 16294 6092 16346
rect 6104 16294 6156 16346
rect 10747 16294 10799 16346
rect 10811 16294 10863 16346
rect 10875 16294 10927 16346
rect 10939 16294 10991 16346
rect 11003 16294 11055 16346
rect 15646 16294 15698 16346
rect 15710 16294 15762 16346
rect 15774 16294 15826 16346
rect 15838 16294 15890 16346
rect 15902 16294 15954 16346
rect 20545 16294 20597 16346
rect 20609 16294 20661 16346
rect 20673 16294 20725 16346
rect 20737 16294 20789 16346
rect 20801 16294 20853 16346
rect 2596 16192 2648 16244
rect 3240 16192 3292 16244
rect 7288 16192 7340 16244
rect 10048 16192 10100 16244
rect 14648 16192 14700 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 20260 16192 20312 16244
rect 3792 16124 3844 16176
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 6828 16056 6880 16108
rect 8668 16167 8720 16176
rect 8668 16133 8677 16167
rect 8677 16133 8711 16167
rect 8711 16133 8720 16167
rect 8668 16124 8720 16133
rect 17776 16124 17828 16176
rect 9772 16056 9824 16108
rect 10508 16056 10560 16108
rect 11612 16056 11664 16108
rect 2504 15988 2556 16040
rect 10416 15988 10468 16040
rect 14280 16056 14332 16108
rect 15108 16056 15160 16108
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 16028 16056 16080 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 17684 16056 17736 16108
rect 19800 16056 19852 16108
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 3399 15750 3451 15802
rect 3463 15750 3515 15802
rect 3527 15750 3579 15802
rect 3591 15750 3643 15802
rect 3655 15750 3707 15802
rect 8298 15750 8350 15802
rect 8362 15750 8414 15802
rect 8426 15750 8478 15802
rect 8490 15750 8542 15802
rect 8554 15750 8606 15802
rect 13197 15750 13249 15802
rect 13261 15750 13313 15802
rect 13325 15750 13377 15802
rect 13389 15750 13441 15802
rect 13453 15750 13505 15802
rect 18096 15750 18148 15802
rect 18160 15750 18212 15802
rect 18224 15750 18276 15802
rect 18288 15750 18340 15802
rect 18352 15750 18404 15802
rect 1952 15648 2004 15700
rect 18696 15648 18748 15700
rect 1492 15444 1544 15496
rect 2688 15444 2740 15496
rect 6828 15444 6880 15496
rect 13728 15580 13780 15632
rect 11612 15512 11664 15564
rect 15108 15555 15160 15564
rect 15108 15521 15117 15555
rect 15117 15521 15151 15555
rect 15151 15521 15160 15555
rect 15108 15512 15160 15521
rect 17040 15580 17092 15632
rect 17592 15512 17644 15564
rect 10508 15444 10560 15496
rect 18512 15444 18564 15496
rect 20076 15487 20128 15496
rect 20076 15453 20085 15487
rect 20085 15453 20119 15487
rect 20119 15453 20128 15487
rect 20076 15444 20128 15453
rect 7288 15376 7340 15428
rect 8116 15376 8168 15428
rect 9772 15376 9824 15428
rect 14096 15376 14148 15428
rect 16120 15376 16172 15428
rect 19340 15376 19392 15428
rect 12348 15351 12400 15360
rect 12348 15317 12357 15351
rect 12357 15317 12391 15351
rect 12391 15317 12400 15351
rect 12348 15308 12400 15317
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 18696 15351 18748 15360
rect 18696 15317 18705 15351
rect 18705 15317 18739 15351
rect 18739 15317 18748 15351
rect 18696 15308 18748 15317
rect 5848 15206 5900 15258
rect 5912 15206 5964 15258
rect 5976 15206 6028 15258
rect 6040 15206 6092 15258
rect 6104 15206 6156 15258
rect 10747 15206 10799 15258
rect 10811 15206 10863 15258
rect 10875 15206 10927 15258
rect 10939 15206 10991 15258
rect 11003 15206 11055 15258
rect 15646 15206 15698 15258
rect 15710 15206 15762 15258
rect 15774 15206 15826 15258
rect 15838 15206 15890 15258
rect 15902 15206 15954 15258
rect 20545 15206 20597 15258
rect 20609 15206 20661 15258
rect 20673 15206 20725 15258
rect 20737 15206 20789 15258
rect 20801 15206 20853 15258
rect 8116 15104 8168 15156
rect 9588 15104 9640 15156
rect 12900 15104 12952 15156
rect 20168 15147 20220 15156
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 5632 15036 5684 15088
rect 18696 15079 18748 15088
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 5356 15011 5408 15020
rect 5356 14977 5365 15011
rect 5365 14977 5399 15011
rect 5399 14977 5408 15011
rect 5356 14968 5408 14977
rect 18696 15045 18705 15079
rect 18705 15045 18739 15079
rect 18739 15045 18748 15079
rect 18696 15036 18748 15045
rect 19340 15036 19392 15088
rect 9128 14900 9180 14952
rect 10876 14968 10928 15020
rect 11152 14968 11204 15020
rect 12348 14968 12400 15020
rect 14096 15011 14148 15020
rect 14096 14977 14114 15011
rect 14114 14977 14148 15011
rect 14096 14968 14148 14977
rect 16488 14900 16540 14952
rect 18420 14943 18472 14952
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 18788 14900 18840 14952
rect 7564 14832 7616 14884
rect 1860 14764 1912 14816
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 7288 14764 7340 14816
rect 9956 14764 10008 14816
rect 11336 14764 11388 14816
rect 12256 14764 12308 14816
rect 14556 14764 14608 14816
rect 3399 14662 3451 14714
rect 3463 14662 3515 14714
rect 3527 14662 3579 14714
rect 3591 14662 3643 14714
rect 3655 14662 3707 14714
rect 8298 14662 8350 14714
rect 8362 14662 8414 14714
rect 8426 14662 8478 14714
rect 8490 14662 8542 14714
rect 8554 14662 8606 14714
rect 13197 14662 13249 14714
rect 13261 14662 13313 14714
rect 13325 14662 13377 14714
rect 13389 14662 13441 14714
rect 13453 14662 13505 14714
rect 18096 14662 18148 14714
rect 18160 14662 18212 14714
rect 18224 14662 18276 14714
rect 18288 14662 18340 14714
rect 18352 14662 18404 14714
rect 10600 14560 10652 14612
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 14096 14560 14148 14612
rect 16580 14560 16632 14612
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 11152 14492 11204 14544
rect 11336 14535 11388 14544
rect 11336 14501 11345 14535
rect 11345 14501 11379 14535
rect 11379 14501 11388 14535
rect 11336 14492 11388 14501
rect 17408 14492 17460 14544
rect 9128 14467 9180 14476
rect 9128 14433 9137 14467
rect 9137 14433 9171 14467
rect 9171 14433 9180 14467
rect 9128 14424 9180 14433
rect 10416 14424 10468 14476
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 17592 14424 17644 14476
rect 1860 14356 1912 14408
rect 7380 14356 7432 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 16856 14356 16908 14408
rect 4528 14288 4580 14340
rect 5356 14288 5408 14340
rect 7288 14288 7340 14340
rect 8760 14288 8812 14340
rect 9864 14288 9916 14340
rect 12532 14288 12584 14340
rect 15200 14288 15252 14340
rect 1952 14220 2004 14272
rect 2872 14220 2924 14272
rect 7196 14220 7248 14272
rect 11520 14220 11572 14272
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 5848 14118 5900 14170
rect 5912 14118 5964 14170
rect 5976 14118 6028 14170
rect 6040 14118 6092 14170
rect 6104 14118 6156 14170
rect 10747 14118 10799 14170
rect 10811 14118 10863 14170
rect 10875 14118 10927 14170
rect 10939 14118 10991 14170
rect 11003 14118 11055 14170
rect 15646 14118 15698 14170
rect 15710 14118 15762 14170
rect 15774 14118 15826 14170
rect 15838 14118 15890 14170
rect 15902 14118 15954 14170
rect 20545 14118 20597 14170
rect 20609 14118 20661 14170
rect 20673 14118 20725 14170
rect 20737 14118 20789 14170
rect 20801 14118 20853 14170
rect 4068 14016 4120 14068
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 5356 14016 5408 14068
rect 7380 14059 7432 14068
rect 7380 14025 7389 14059
rect 7389 14025 7423 14059
rect 7423 14025 7432 14059
rect 7380 14016 7432 14025
rect 10416 14016 10468 14068
rect 14372 14016 14424 14068
rect 3792 13948 3844 14000
rect 9864 13948 9916 14000
rect 14648 13948 14700 14000
rect 18420 13948 18472 14000
rect 19340 13948 19392 14000
rect 1492 13880 1544 13932
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 6828 13880 6880 13932
rect 7196 13923 7248 13932
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 8208 13880 8260 13932
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 11060 13880 11112 13932
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 6460 13812 6512 13864
rect 8116 13812 8168 13864
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 12440 13812 12492 13864
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 18788 13812 18840 13864
rect 20168 13719 20220 13728
rect 20168 13685 20177 13719
rect 20177 13685 20211 13719
rect 20211 13685 20220 13719
rect 20168 13676 20220 13685
rect 3399 13574 3451 13626
rect 3463 13574 3515 13626
rect 3527 13574 3579 13626
rect 3591 13574 3643 13626
rect 3655 13574 3707 13626
rect 8298 13574 8350 13626
rect 8362 13574 8414 13626
rect 8426 13574 8478 13626
rect 8490 13574 8542 13626
rect 8554 13574 8606 13626
rect 13197 13574 13249 13626
rect 13261 13574 13313 13626
rect 13325 13574 13377 13626
rect 13389 13574 13441 13626
rect 13453 13574 13505 13626
rect 18096 13574 18148 13626
rect 18160 13574 18212 13626
rect 18224 13574 18276 13626
rect 18288 13574 18340 13626
rect 18352 13574 18404 13626
rect 4712 13472 4764 13524
rect 11060 13515 11112 13524
rect 11060 13481 11069 13515
rect 11069 13481 11103 13515
rect 11103 13481 11112 13515
rect 11060 13472 11112 13481
rect 12808 13472 12860 13524
rect 13452 13472 13504 13524
rect 14096 13472 14148 13524
rect 19984 13515 20036 13524
rect 1492 13404 1544 13456
rect 10600 13404 10652 13456
rect 12440 13447 12492 13456
rect 12440 13413 12449 13447
rect 12449 13413 12483 13447
rect 12483 13413 12492 13447
rect 12440 13404 12492 13413
rect 5540 13379 5592 13388
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 7196 13336 7248 13388
rect 10416 13336 10468 13388
rect 15200 13336 15252 13388
rect 19984 13481 19993 13515
rect 19993 13481 20027 13515
rect 20027 13481 20036 13515
rect 19984 13472 20036 13481
rect 1952 13311 2004 13320
rect 1952 13277 1961 13311
rect 1961 13277 1995 13311
rect 1995 13277 2004 13311
rect 1952 13268 2004 13277
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 4528 13268 4580 13320
rect 7288 13268 7340 13320
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 13084 13268 13136 13320
rect 13452 13311 13504 13320
rect 13452 13277 13460 13311
rect 13460 13277 13504 13311
rect 13452 13268 13504 13277
rect 13912 13268 13964 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 20168 13311 20220 13320
rect 20168 13277 20177 13311
rect 20177 13277 20211 13311
rect 20211 13277 20220 13311
rect 20168 13268 20220 13277
rect 7748 13200 7800 13252
rect 15200 13200 15252 13252
rect 16120 13200 16172 13252
rect 7104 13132 7156 13184
rect 16672 13132 16724 13184
rect 18604 13132 18656 13184
rect 5848 13030 5900 13082
rect 5912 13030 5964 13082
rect 5976 13030 6028 13082
rect 6040 13030 6092 13082
rect 6104 13030 6156 13082
rect 10747 13030 10799 13082
rect 10811 13030 10863 13082
rect 10875 13030 10927 13082
rect 10939 13030 10991 13082
rect 11003 13030 11055 13082
rect 15646 13030 15698 13082
rect 15710 13030 15762 13082
rect 15774 13030 15826 13082
rect 15838 13030 15890 13082
rect 15902 13030 15954 13082
rect 20545 13030 20597 13082
rect 20609 13030 20661 13082
rect 20673 13030 20725 13082
rect 20737 13030 20789 13082
rect 20801 13030 20853 13082
rect 2044 12792 2096 12844
rect 14648 12928 14700 12980
rect 7104 12860 7156 12912
rect 7564 12860 7616 12912
rect 14096 12860 14148 12912
rect 16948 12928 17000 12980
rect 19340 12860 19392 12912
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9956 12835 10008 12844
rect 9956 12801 9965 12835
rect 9965 12801 9999 12835
rect 9999 12801 10008 12835
rect 9956 12792 10008 12801
rect 15568 12792 15620 12844
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 11244 12724 11296 12776
rect 12624 12724 12676 12776
rect 16120 12724 16172 12776
rect 17776 12724 17828 12776
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 18696 12767 18748 12776
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 11704 12699 11756 12708
rect 11704 12665 11713 12699
rect 11713 12665 11747 12699
rect 11747 12665 11756 12699
rect 11704 12656 11756 12665
rect 1584 12588 1636 12640
rect 5172 12588 5224 12640
rect 8668 12588 8720 12640
rect 9128 12588 9180 12640
rect 9956 12588 10008 12640
rect 10508 12588 10560 12640
rect 20168 12631 20220 12640
rect 20168 12597 20177 12631
rect 20177 12597 20211 12631
rect 20211 12597 20220 12631
rect 20168 12588 20220 12597
rect 3399 12486 3451 12538
rect 3463 12486 3515 12538
rect 3527 12486 3579 12538
rect 3591 12486 3643 12538
rect 3655 12486 3707 12538
rect 8298 12486 8350 12538
rect 8362 12486 8414 12538
rect 8426 12486 8478 12538
rect 8490 12486 8542 12538
rect 8554 12486 8606 12538
rect 13197 12486 13249 12538
rect 13261 12486 13313 12538
rect 13325 12486 13377 12538
rect 13389 12486 13441 12538
rect 13453 12486 13505 12538
rect 18096 12486 18148 12538
rect 18160 12486 18212 12538
rect 18224 12486 18276 12538
rect 18288 12486 18340 12538
rect 18352 12486 18404 12538
rect 6552 12384 6604 12436
rect 8760 12384 8812 12436
rect 11152 12384 11204 12436
rect 11704 12384 11756 12436
rect 14188 12384 14240 12436
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 18696 12384 18748 12436
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 13084 12316 13136 12368
rect 9956 12248 10008 12300
rect 18144 12316 18196 12368
rect 19984 12359 20036 12368
rect 19984 12325 19993 12359
rect 19993 12325 20027 12359
rect 20027 12325 20036 12359
rect 19984 12316 20036 12325
rect 18052 12248 18104 12300
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 4804 12180 4856 12232
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 6184 12180 6236 12232
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 3516 12044 3568 12096
rect 5264 12044 5316 12096
rect 6828 12180 6880 12232
rect 7104 12180 7156 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 18604 12180 18656 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 9864 12112 9916 12164
rect 11980 12155 12032 12164
rect 11980 12121 11989 12155
rect 11989 12121 12023 12155
rect 12023 12121 12032 12155
rect 11980 12112 12032 12121
rect 12624 12112 12676 12164
rect 14004 12112 14056 12164
rect 14096 12044 14148 12096
rect 16120 12112 16172 12164
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 5848 11942 5900 11994
rect 5912 11942 5964 11994
rect 5976 11942 6028 11994
rect 6040 11942 6092 11994
rect 6104 11942 6156 11994
rect 10747 11942 10799 11994
rect 10811 11942 10863 11994
rect 10875 11942 10927 11994
rect 10939 11942 10991 11994
rect 11003 11942 11055 11994
rect 15646 11942 15698 11994
rect 15710 11942 15762 11994
rect 15774 11942 15826 11994
rect 15838 11942 15890 11994
rect 15902 11942 15954 11994
rect 20545 11942 20597 11994
rect 20609 11942 20661 11994
rect 20673 11942 20725 11994
rect 20737 11942 20789 11994
rect 20801 11942 20853 11994
rect 4344 11840 4396 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 6828 11840 6880 11892
rect 11244 11840 11296 11892
rect 11980 11840 12032 11892
rect 18144 11840 18196 11892
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 4620 11704 4672 11756
rect 6184 11704 6236 11756
rect 6828 11704 6880 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 13084 11704 13136 11756
rect 13912 11772 13964 11824
rect 11152 11636 11204 11688
rect 11704 11636 11756 11688
rect 15016 11704 15068 11756
rect 16580 11704 16632 11756
rect 16948 11704 17000 11756
rect 14004 11636 14056 11688
rect 8208 11568 8260 11620
rect 6184 11500 6236 11552
rect 10416 11500 10468 11552
rect 16856 11636 16908 11688
rect 18052 11636 18104 11688
rect 15844 11568 15896 11620
rect 18696 11500 18748 11552
rect 3399 11398 3451 11450
rect 3463 11398 3515 11450
rect 3527 11398 3579 11450
rect 3591 11398 3643 11450
rect 3655 11398 3707 11450
rect 8298 11398 8350 11450
rect 8362 11398 8414 11450
rect 8426 11398 8478 11450
rect 8490 11398 8542 11450
rect 8554 11398 8606 11450
rect 13197 11398 13249 11450
rect 13261 11398 13313 11450
rect 13325 11398 13377 11450
rect 13389 11398 13441 11450
rect 13453 11398 13505 11450
rect 18096 11398 18148 11450
rect 18160 11398 18212 11450
rect 18224 11398 18276 11450
rect 18288 11398 18340 11450
rect 18352 11398 18404 11450
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 6828 11296 6880 11348
rect 15016 11296 15068 11348
rect 15844 11339 15896 11348
rect 15844 11305 15853 11339
rect 15853 11305 15887 11339
rect 15887 11305 15896 11339
rect 15844 11296 15896 11305
rect 17776 11296 17828 11348
rect 1492 11228 1544 11280
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 16212 11228 16264 11280
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 8116 11160 8168 11212
rect 11244 11160 11296 11212
rect 16948 11160 17000 11212
rect 17960 11160 18012 11212
rect 8668 11092 8720 11144
rect 11428 11135 11480 11144
rect 11428 11101 11446 11135
rect 11446 11101 11480 11135
rect 11428 11092 11480 11101
rect 16028 11092 16080 11144
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 7748 11024 7800 11076
rect 9496 11024 9548 11076
rect 9864 11024 9916 11076
rect 10232 11024 10284 11076
rect 15200 11024 15252 11076
rect 15568 11024 15620 11076
rect 8668 10956 8720 11008
rect 11888 10956 11940 11008
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 5848 10854 5900 10906
rect 5912 10854 5964 10906
rect 5976 10854 6028 10906
rect 6040 10854 6092 10906
rect 6104 10854 6156 10906
rect 10747 10854 10799 10906
rect 10811 10854 10863 10906
rect 10875 10854 10927 10906
rect 10939 10854 10991 10906
rect 11003 10854 11055 10906
rect 15646 10854 15698 10906
rect 15710 10854 15762 10906
rect 15774 10854 15826 10906
rect 15838 10854 15890 10906
rect 15902 10854 15954 10906
rect 20545 10854 20597 10906
rect 20609 10854 20661 10906
rect 20673 10854 20725 10906
rect 20737 10854 20789 10906
rect 20801 10854 20853 10906
rect 3976 10795 4028 10804
rect 3976 10761 3985 10795
rect 3985 10761 4019 10795
rect 4019 10761 4028 10795
rect 3976 10752 4028 10761
rect 17868 10752 17920 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2320 10616 2372 10668
rect 3240 10616 3292 10668
rect 8208 10616 8260 10668
rect 8760 10684 8812 10736
rect 7380 10548 7432 10600
rect 9220 10548 9272 10600
rect 12624 10684 12676 10736
rect 14648 10684 14700 10736
rect 18696 10727 18748 10736
rect 18696 10693 18705 10727
rect 18705 10693 18739 10727
rect 18739 10693 18748 10727
rect 18696 10684 18748 10693
rect 19340 10684 19392 10736
rect 11612 10616 11664 10668
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 18788 10548 18840 10600
rect 1952 10412 2004 10464
rect 2780 10412 2832 10464
rect 9588 10412 9640 10464
rect 14280 10412 14332 10464
rect 15568 10412 15620 10464
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 3399 10310 3451 10362
rect 3463 10310 3515 10362
rect 3527 10310 3579 10362
rect 3591 10310 3643 10362
rect 3655 10310 3707 10362
rect 8298 10310 8350 10362
rect 8362 10310 8414 10362
rect 8426 10310 8478 10362
rect 8490 10310 8542 10362
rect 8554 10310 8606 10362
rect 13197 10310 13249 10362
rect 13261 10310 13313 10362
rect 13325 10310 13377 10362
rect 13389 10310 13441 10362
rect 13453 10310 13505 10362
rect 18096 10310 18148 10362
rect 18160 10310 18212 10362
rect 18224 10310 18276 10362
rect 18288 10310 18340 10362
rect 18352 10310 18404 10362
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 3240 10208 3292 10260
rect 11428 10251 11480 10260
rect 11428 10217 11437 10251
rect 11437 10217 11471 10251
rect 11471 10217 11480 10251
rect 11428 10208 11480 10217
rect 12624 10208 12676 10260
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 11888 10183 11940 10192
rect 11888 10149 11897 10183
rect 11897 10149 11931 10183
rect 11931 10149 11940 10183
rect 11888 10140 11940 10149
rect 11612 10072 11664 10124
rect 15200 10072 15252 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 8668 10004 8720 10056
rect 9588 10004 9640 10056
rect 9956 10047 10008 10056
rect 9956 10013 9965 10047
rect 9965 10013 9999 10047
rect 9999 10013 10008 10047
rect 9956 10004 10008 10013
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 20168 10047 20220 10056
rect 20168 10013 20177 10047
rect 20177 10013 20211 10047
rect 20211 10013 20220 10047
rect 20168 10004 20220 10013
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 15200 9936 15252 9988
rect 8760 9868 8812 9920
rect 9312 9868 9364 9920
rect 10508 9868 10560 9920
rect 11980 9868 12032 9920
rect 5848 9766 5900 9818
rect 5912 9766 5964 9818
rect 5976 9766 6028 9818
rect 6040 9766 6092 9818
rect 6104 9766 6156 9818
rect 10747 9766 10799 9818
rect 10811 9766 10863 9818
rect 10875 9766 10927 9818
rect 10939 9766 10991 9818
rect 11003 9766 11055 9818
rect 15646 9766 15698 9818
rect 15710 9766 15762 9818
rect 15774 9766 15826 9818
rect 15838 9766 15890 9818
rect 15902 9766 15954 9818
rect 20545 9766 20597 9818
rect 20609 9766 20661 9818
rect 20673 9766 20725 9818
rect 20737 9766 20789 9818
rect 20801 9766 20853 9818
rect 9956 9707 10008 9716
rect 9956 9673 9965 9707
rect 9965 9673 9999 9707
rect 9999 9673 10008 9707
rect 9956 9664 10008 9673
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 1860 9528 1912 9580
rect 4896 9596 4948 9648
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 10508 9596 10560 9648
rect 5540 9528 5592 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 17224 9596 17276 9648
rect 19340 9596 19392 9648
rect 17960 9571 18012 9580
rect 17960 9537 17969 9571
rect 17969 9537 18003 9571
rect 18003 9537 18012 9571
rect 17960 9528 18012 9537
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 3240 9460 3292 9512
rect 4528 9460 4580 9512
rect 11980 9460 12032 9512
rect 17868 9460 17920 9512
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 7288 9324 7340 9376
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 3399 9222 3451 9274
rect 3463 9222 3515 9274
rect 3527 9222 3579 9274
rect 3591 9222 3643 9274
rect 3655 9222 3707 9274
rect 8298 9222 8350 9274
rect 8362 9222 8414 9274
rect 8426 9222 8478 9274
rect 8490 9222 8542 9274
rect 8554 9222 8606 9274
rect 13197 9222 13249 9274
rect 13261 9222 13313 9274
rect 13325 9222 13377 9274
rect 13389 9222 13441 9274
rect 13453 9222 13505 9274
rect 18096 9222 18148 9274
rect 18160 9222 18212 9274
rect 18224 9222 18276 9274
rect 18288 9222 18340 9274
rect 18352 9222 18404 9274
rect 3240 9120 3292 9172
rect 7472 9120 7524 9172
rect 17960 9120 18012 9172
rect 13820 9052 13872 9104
rect 17868 9052 17920 9104
rect 3148 8984 3200 9036
rect 9588 8984 9640 9036
rect 12256 8984 12308 9036
rect 16028 8984 16080 9036
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 10324 8916 10376 8968
rect 12072 8916 12124 8968
rect 13544 8916 13596 8968
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 17132 8916 17184 8968
rect 18420 8959 18472 8968
rect 5264 8848 5316 8900
rect 5448 8848 5500 8900
rect 6920 8848 6972 8900
rect 9956 8848 10008 8900
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 9772 8780 9824 8832
rect 12808 8780 12860 8832
rect 16120 8780 16172 8832
rect 17592 8848 17644 8900
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 19340 8848 19392 8900
rect 19616 8891 19668 8900
rect 19616 8857 19625 8891
rect 19625 8857 19659 8891
rect 19659 8857 19668 8891
rect 19616 8848 19668 8857
rect 19248 8780 19300 8832
rect 5848 8678 5900 8730
rect 5912 8678 5964 8730
rect 5976 8678 6028 8730
rect 6040 8678 6092 8730
rect 6104 8678 6156 8730
rect 10747 8678 10799 8730
rect 10811 8678 10863 8730
rect 10875 8678 10927 8730
rect 10939 8678 10991 8730
rect 11003 8678 11055 8730
rect 15646 8678 15698 8730
rect 15710 8678 15762 8730
rect 15774 8678 15826 8730
rect 15838 8678 15890 8730
rect 15902 8678 15954 8730
rect 20545 8678 20597 8730
rect 20609 8678 20661 8730
rect 20673 8678 20725 8730
rect 20737 8678 20789 8730
rect 20801 8678 20853 8730
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 2780 8576 2832 8628
rect 5264 8576 5316 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 12072 8619 12124 8628
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 15108 8576 15160 8628
rect 19984 8619 20036 8628
rect 19984 8585 19993 8619
rect 19993 8585 20027 8619
rect 20027 8585 20036 8619
rect 19984 8576 20036 8585
rect 4804 8508 4856 8560
rect 7932 8508 7984 8560
rect 8668 8508 8720 8560
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 9496 8440 9548 8492
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 12808 8508 12860 8560
rect 15660 8508 15712 8560
rect 16120 8508 16172 8560
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 17592 8508 17644 8560
rect 3148 8372 3200 8424
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 2872 8347 2924 8356
rect 2872 8313 2881 8347
rect 2881 8313 2915 8347
rect 2915 8313 2924 8347
rect 2872 8304 2924 8313
rect 5356 8304 5408 8356
rect 12440 8372 12492 8424
rect 12900 8372 12952 8424
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 20168 8483 20220 8492
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 9680 8236 9732 8288
rect 10508 8279 10560 8288
rect 10508 8245 10517 8279
rect 10517 8245 10551 8279
rect 10551 8245 10560 8279
rect 10508 8236 10560 8245
rect 14556 8236 14608 8288
rect 17776 8236 17828 8288
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 3399 8134 3451 8186
rect 3463 8134 3515 8186
rect 3527 8134 3579 8186
rect 3591 8134 3643 8186
rect 3655 8134 3707 8186
rect 8298 8134 8350 8186
rect 8362 8134 8414 8186
rect 8426 8134 8478 8186
rect 8490 8134 8542 8186
rect 8554 8134 8606 8186
rect 13197 8134 13249 8186
rect 13261 8134 13313 8186
rect 13325 8134 13377 8186
rect 13389 8134 13441 8186
rect 13453 8134 13505 8186
rect 18096 8134 18148 8186
rect 18160 8134 18212 8186
rect 18224 8134 18276 8186
rect 18288 8134 18340 8186
rect 18352 8134 18404 8186
rect 4252 8032 4304 8084
rect 7564 8032 7616 8084
rect 3240 7964 3292 8016
rect 5448 7896 5500 7948
rect 8116 7896 8168 7948
rect 8668 8032 8720 8084
rect 10324 8032 10376 8084
rect 11152 8032 11204 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 13544 8032 13596 8084
rect 16028 8075 16080 8084
rect 16028 8041 16037 8075
rect 16037 8041 16071 8075
rect 16071 8041 16080 8075
rect 16028 8032 16080 8041
rect 18512 8032 18564 8084
rect 19616 8032 19668 8084
rect 1676 7828 1728 7880
rect 3148 7828 3200 7880
rect 4344 7871 4396 7880
rect 4344 7837 4352 7871
rect 4352 7837 4396 7871
rect 4344 7828 4396 7837
rect 5632 7828 5684 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 9496 7760 9548 7812
rect 9956 7964 10008 8016
rect 10508 7896 10560 7948
rect 18420 8007 18472 8016
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 15660 7828 15712 7880
rect 16028 7828 16080 7880
rect 18420 7973 18429 8007
rect 18429 7973 18463 8007
rect 18463 7973 18472 8007
rect 18420 7964 18472 7973
rect 19064 7828 19116 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 2320 7692 2372 7744
rect 3976 7692 4028 7744
rect 5848 7590 5900 7642
rect 5912 7590 5964 7642
rect 5976 7590 6028 7642
rect 6040 7590 6092 7642
rect 6104 7590 6156 7642
rect 10747 7590 10799 7642
rect 10811 7590 10863 7642
rect 10875 7590 10927 7642
rect 10939 7590 10991 7642
rect 11003 7590 11055 7642
rect 15646 7590 15698 7642
rect 15710 7590 15762 7642
rect 15774 7590 15826 7642
rect 15838 7590 15890 7642
rect 15902 7590 15954 7642
rect 20545 7590 20597 7642
rect 20609 7590 20661 7642
rect 20673 7590 20725 7642
rect 20737 7590 20789 7642
rect 20801 7590 20853 7642
rect 6828 7488 6880 7540
rect 9496 7488 9548 7540
rect 11152 7531 11204 7540
rect 2504 7420 2556 7472
rect 9680 7463 9732 7472
rect 9680 7429 9689 7463
rect 9689 7429 9723 7463
rect 9723 7429 9732 7463
rect 9680 7420 9732 7429
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 19616 7488 19668 7540
rect 5632 7352 5684 7404
rect 7288 7352 7340 7404
rect 7472 7352 7524 7404
rect 8668 7352 8720 7404
rect 19340 7420 19392 7472
rect 14556 7352 14608 7404
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 5540 7284 5592 7336
rect 5724 7284 5776 7336
rect 9772 7284 9824 7336
rect 17132 7284 17184 7336
rect 17868 7284 17920 7336
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 4344 7259 4396 7268
rect 4344 7225 4353 7259
rect 4353 7225 4387 7259
rect 4387 7225 4396 7259
rect 4344 7216 4396 7225
rect 1676 7148 1728 7200
rect 3240 7148 3292 7200
rect 3792 7148 3844 7200
rect 4804 7148 4856 7200
rect 5632 7148 5684 7200
rect 9128 7148 9180 7200
rect 11428 7148 11480 7200
rect 15660 7148 15712 7200
rect 20168 7191 20220 7200
rect 20168 7157 20177 7191
rect 20177 7157 20211 7191
rect 20211 7157 20220 7191
rect 20168 7148 20220 7157
rect 3399 7046 3451 7098
rect 3463 7046 3515 7098
rect 3527 7046 3579 7098
rect 3591 7046 3643 7098
rect 3655 7046 3707 7098
rect 8298 7046 8350 7098
rect 8362 7046 8414 7098
rect 8426 7046 8478 7098
rect 8490 7046 8542 7098
rect 8554 7046 8606 7098
rect 13197 7046 13249 7098
rect 13261 7046 13313 7098
rect 13325 7046 13377 7098
rect 13389 7046 13441 7098
rect 13453 7046 13505 7098
rect 18096 7046 18148 7098
rect 18160 7046 18212 7098
rect 18224 7046 18276 7098
rect 18288 7046 18340 7098
rect 18352 7046 18404 7098
rect 3148 6944 3200 6996
rect 4344 6944 4396 6996
rect 1676 6876 1728 6928
rect 12348 6944 12400 6996
rect 12256 6876 12308 6928
rect 13820 6876 13872 6928
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 5724 6808 5776 6860
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 3976 6783 4028 6792
rect 3976 6749 4020 6783
rect 4020 6749 4028 6783
rect 5356 6783 5408 6792
rect 3976 6740 4028 6749
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 9220 6808 9272 6860
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9680 6740 9732 6792
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 7472 6672 7524 6724
rect 15292 6672 15344 6724
rect 7932 6604 7984 6656
rect 10600 6604 10652 6656
rect 16856 6604 16908 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 5848 6502 5900 6554
rect 5912 6502 5964 6554
rect 5976 6502 6028 6554
rect 6040 6502 6092 6554
rect 6104 6502 6156 6554
rect 10747 6502 10799 6554
rect 10811 6502 10863 6554
rect 10875 6502 10927 6554
rect 10939 6502 10991 6554
rect 11003 6502 11055 6554
rect 15646 6502 15698 6554
rect 15710 6502 15762 6554
rect 15774 6502 15826 6554
rect 15838 6502 15890 6554
rect 15902 6502 15954 6554
rect 20545 6502 20597 6554
rect 20609 6502 20661 6554
rect 20673 6502 20725 6554
rect 20737 6502 20789 6554
rect 20801 6502 20853 6554
rect 2872 6400 2924 6452
rect 7472 6400 7524 6452
rect 15384 6400 15436 6452
rect 18696 6400 18748 6452
rect 2872 6264 2924 6316
rect 3240 6264 3292 6316
rect 10508 6332 10560 6384
rect 12532 6332 12584 6384
rect 16580 6332 16632 6384
rect 17040 6332 17092 6384
rect 3976 6264 4028 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 13912 6264 13964 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 3148 6196 3200 6248
rect 3792 6196 3844 6248
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 14188 6196 14240 6248
rect 15292 6196 15344 6248
rect 5080 6171 5132 6180
rect 5080 6137 5089 6171
rect 5089 6137 5123 6171
rect 5123 6137 5132 6171
rect 5080 6128 5132 6137
rect 9772 6171 9824 6180
rect 9772 6137 9781 6171
rect 9781 6137 9815 6171
rect 9815 6137 9824 6171
rect 9772 6128 9824 6137
rect 15016 6128 15068 6180
rect 16120 6128 16172 6180
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 5632 6060 5684 6112
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8760 6060 8812 6112
rect 9680 6060 9732 6112
rect 10508 6060 10560 6112
rect 16212 6060 16264 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 3399 5958 3451 6010
rect 3463 5958 3515 6010
rect 3527 5958 3579 6010
rect 3591 5958 3643 6010
rect 3655 5958 3707 6010
rect 8298 5958 8350 6010
rect 8362 5958 8414 6010
rect 8426 5958 8478 6010
rect 8490 5958 8542 6010
rect 8554 5958 8606 6010
rect 13197 5958 13249 6010
rect 13261 5958 13313 6010
rect 13325 5958 13377 6010
rect 13389 5958 13441 6010
rect 13453 5958 13505 6010
rect 18096 5958 18148 6010
rect 18160 5958 18212 6010
rect 18224 5958 18276 6010
rect 18288 5958 18340 6010
rect 18352 5958 18404 6010
rect 6460 5856 6512 5908
rect 9956 5856 10008 5908
rect 13912 5856 13964 5908
rect 15016 5899 15068 5908
rect 15016 5865 15025 5899
rect 15025 5865 15059 5899
rect 15059 5865 15068 5899
rect 15016 5856 15068 5865
rect 5264 5788 5316 5840
rect 3148 5763 3200 5772
rect 3148 5729 3157 5763
rect 3157 5729 3191 5763
rect 3191 5729 3200 5763
rect 3148 5720 3200 5729
rect 6184 5763 6236 5772
rect 6184 5729 6193 5763
rect 6193 5729 6227 5763
rect 6227 5729 6236 5763
rect 6184 5720 6236 5729
rect 7932 5788 7984 5840
rect 16028 5831 16080 5840
rect 9772 5720 9824 5772
rect 16028 5797 16037 5831
rect 16037 5797 16071 5831
rect 16071 5797 16080 5831
rect 16028 5788 16080 5797
rect 15292 5720 15344 5772
rect 18604 5720 18656 5772
rect 2872 5652 2924 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4712 5584 4764 5636
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 13912 5652 13964 5704
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 9404 5584 9456 5636
rect 10600 5584 10652 5636
rect 12440 5584 12492 5636
rect 19340 5584 19392 5636
rect 5080 5516 5132 5568
rect 17500 5516 17552 5568
rect 18880 5559 18932 5568
rect 18880 5525 18889 5559
rect 18889 5525 18923 5559
rect 18923 5525 18932 5559
rect 18880 5516 18932 5525
rect 5848 5414 5900 5466
rect 5912 5414 5964 5466
rect 5976 5414 6028 5466
rect 6040 5414 6092 5466
rect 6104 5414 6156 5466
rect 10747 5414 10799 5466
rect 10811 5414 10863 5466
rect 10875 5414 10927 5466
rect 10939 5414 10991 5466
rect 11003 5414 11055 5466
rect 15646 5414 15698 5466
rect 15710 5414 15762 5466
rect 15774 5414 15826 5466
rect 15838 5414 15890 5466
rect 15902 5414 15954 5466
rect 20545 5414 20597 5466
rect 20609 5414 20661 5466
rect 20673 5414 20725 5466
rect 20737 5414 20789 5466
rect 20801 5414 20853 5466
rect 2504 5312 2556 5364
rect 4712 5312 4764 5364
rect 5264 5312 5316 5364
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 5632 5219 5684 5228
rect 7840 5244 7892 5296
rect 8760 5312 8812 5364
rect 9404 5355 9456 5364
rect 9404 5321 9413 5355
rect 9413 5321 9447 5355
rect 9447 5321 9456 5355
rect 9404 5312 9456 5321
rect 12440 5244 12492 5296
rect 13912 5312 13964 5364
rect 16948 5244 17000 5296
rect 17500 5287 17552 5296
rect 17500 5253 17509 5287
rect 17509 5253 17543 5287
rect 17543 5253 17552 5287
rect 17500 5244 17552 5253
rect 19340 5244 19392 5296
rect 5632 5185 5676 5219
rect 5676 5185 5684 5219
rect 5632 5176 5684 5185
rect 9956 5176 10008 5228
rect 10508 5176 10560 5228
rect 13820 5176 13872 5228
rect 17132 5176 17184 5228
rect 7932 5108 7984 5160
rect 9404 5108 9456 5160
rect 10600 5108 10652 5160
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 16120 5108 16172 5160
rect 10232 5015 10284 5024
rect 10232 4981 10241 5015
rect 10241 4981 10275 5015
rect 10275 4981 10284 5015
rect 10232 4972 10284 4981
rect 15936 4972 15988 5024
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 3399 4870 3451 4922
rect 3463 4870 3515 4922
rect 3527 4870 3579 4922
rect 3591 4870 3643 4922
rect 3655 4870 3707 4922
rect 8298 4870 8350 4922
rect 8362 4870 8414 4922
rect 8426 4870 8478 4922
rect 8490 4870 8542 4922
rect 8554 4870 8606 4922
rect 13197 4870 13249 4922
rect 13261 4870 13313 4922
rect 13325 4870 13377 4922
rect 13389 4870 13441 4922
rect 13453 4870 13505 4922
rect 18096 4870 18148 4922
rect 18160 4870 18212 4922
rect 18224 4870 18276 4922
rect 18288 4870 18340 4922
rect 18352 4870 18404 4922
rect 6184 4768 6236 4820
rect 8944 4768 8996 4820
rect 16028 4768 16080 4820
rect 15936 4743 15988 4752
rect 15936 4709 15945 4743
rect 15945 4709 15979 4743
rect 15979 4709 15988 4743
rect 15936 4700 15988 4709
rect 2780 4632 2832 4684
rect 8760 4632 8812 4684
rect 15200 4632 15252 4684
rect 3148 4564 3200 4616
rect 5080 4564 5132 4616
rect 5448 4564 5500 4616
rect 10232 4564 10284 4616
rect 15384 4564 15436 4616
rect 2504 4496 2556 4548
rect 6644 4539 6696 4548
rect 6644 4505 6653 4539
rect 6653 4505 6687 4539
rect 6687 4505 6696 4539
rect 6644 4496 6696 4505
rect 7932 4496 7984 4548
rect 1676 4428 1728 4480
rect 17684 4428 17736 4480
rect 5848 4326 5900 4378
rect 5912 4326 5964 4378
rect 5976 4326 6028 4378
rect 6040 4326 6092 4378
rect 6104 4326 6156 4378
rect 10747 4326 10799 4378
rect 10811 4326 10863 4378
rect 10875 4326 10927 4378
rect 10939 4326 10991 4378
rect 11003 4326 11055 4378
rect 15646 4326 15698 4378
rect 15710 4326 15762 4378
rect 15774 4326 15826 4378
rect 15838 4326 15890 4378
rect 15902 4326 15954 4378
rect 20545 4326 20597 4378
rect 20609 4326 20661 4378
rect 20673 4326 20725 4378
rect 20737 4326 20789 4378
rect 20801 4326 20853 4378
rect 6644 4224 6696 4276
rect 2504 4156 2556 4208
rect 8760 4156 8812 4208
rect 19340 4156 19392 4208
rect 3148 4088 3200 4140
rect 6460 4088 6512 4140
rect 7380 4020 7432 4072
rect 8208 4020 8260 4072
rect 17132 4088 17184 4140
rect 10416 4020 10468 4072
rect 17684 3952 17736 4004
rect 2320 3884 2372 3936
rect 2964 3884 3016 3936
rect 9680 3884 9732 3936
rect 9956 3884 10008 3936
rect 19892 3884 19944 3936
rect 3399 3782 3451 3834
rect 3463 3782 3515 3834
rect 3527 3782 3579 3834
rect 3591 3782 3643 3834
rect 3655 3782 3707 3834
rect 8298 3782 8350 3834
rect 8362 3782 8414 3834
rect 8426 3782 8478 3834
rect 8490 3782 8542 3834
rect 8554 3782 8606 3834
rect 13197 3782 13249 3834
rect 13261 3782 13313 3834
rect 13325 3782 13377 3834
rect 13389 3782 13441 3834
rect 13453 3782 13505 3834
rect 18096 3782 18148 3834
rect 18160 3782 18212 3834
rect 18224 3782 18276 3834
rect 18288 3782 18340 3834
rect 18352 3782 18404 3834
rect 572 3612 624 3664
rect 10600 3612 10652 3664
rect 4252 3544 4304 3596
rect 5448 3544 5500 3596
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 3240 3476 3292 3528
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 11520 3544 11572 3596
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 16028 3544 16080 3596
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 5356 3451 5408 3460
rect 5356 3417 5365 3451
rect 5365 3417 5399 3451
rect 5399 3417 5408 3451
rect 5356 3408 5408 3417
rect 6920 3408 6972 3460
rect 11336 3408 11388 3460
rect 16856 3408 16908 3460
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 7104 3340 7156 3392
rect 12532 3340 12584 3392
rect 17408 3340 17460 3392
rect 20076 3383 20128 3392
rect 20076 3349 20085 3383
rect 20085 3349 20119 3383
rect 20119 3349 20128 3383
rect 20076 3340 20128 3349
rect 5848 3238 5900 3290
rect 5912 3238 5964 3290
rect 5976 3238 6028 3290
rect 6040 3238 6092 3290
rect 6104 3238 6156 3290
rect 10747 3238 10799 3290
rect 10811 3238 10863 3290
rect 10875 3238 10927 3290
rect 10939 3238 10991 3290
rect 11003 3238 11055 3290
rect 15646 3238 15698 3290
rect 15710 3238 15762 3290
rect 15774 3238 15826 3290
rect 15838 3238 15890 3290
rect 15902 3238 15954 3290
rect 20545 3238 20597 3290
rect 20609 3238 20661 3290
rect 20673 3238 20725 3290
rect 20737 3238 20789 3290
rect 20801 3238 20853 3290
rect 2504 3136 2556 3188
rect 4620 3136 4672 3188
rect 16856 3136 16908 3188
rect 5356 3068 5408 3120
rect 11336 3068 11388 3120
rect 12440 3068 12492 3120
rect 1676 3000 1728 3052
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2964 3000 3016 3052
rect 3148 3000 3200 3052
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 7932 3000 7984 3052
rect 9772 3000 9824 3052
rect 16764 3000 16816 3052
rect 18880 3000 18932 3052
rect 19800 3000 19852 3052
rect 3792 2932 3844 2984
rect 4252 2932 4304 2984
rect 8208 2932 8260 2984
rect 16028 2932 16080 2984
rect 19432 2932 19484 2984
rect 19248 2864 19300 2916
rect 21180 2864 21232 2916
rect 1860 2796 1912 2848
rect 3056 2796 3108 2848
rect 5724 2796 5776 2848
rect 8668 2796 8720 2848
rect 11152 2796 11204 2848
rect 19156 2796 19208 2848
rect 19892 2796 19944 2848
rect 3399 2694 3451 2746
rect 3463 2694 3515 2746
rect 3527 2694 3579 2746
rect 3591 2694 3643 2746
rect 3655 2694 3707 2746
rect 8298 2694 8350 2746
rect 8362 2694 8414 2746
rect 8426 2694 8478 2746
rect 8490 2694 8542 2746
rect 8554 2694 8606 2746
rect 13197 2694 13249 2746
rect 13261 2694 13313 2746
rect 13325 2694 13377 2746
rect 13389 2694 13441 2746
rect 13453 2694 13505 2746
rect 18096 2694 18148 2746
rect 18160 2694 18212 2746
rect 18224 2694 18276 2746
rect 18288 2694 18340 2746
rect 18352 2694 18404 2746
rect 3240 2592 3292 2644
rect 3792 2592 3844 2644
rect 5356 2592 5408 2644
rect 6000 2592 6052 2644
rect 19248 2592 19300 2644
rect 9496 2456 9548 2508
rect 7104 2431 7156 2440
rect 2504 2320 2556 2372
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 8668 2388 8720 2440
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 15384 2388 15436 2440
rect 16672 2388 16724 2440
rect 17408 2388 17460 2440
rect 19708 2456 19760 2508
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 4252 2320 4304 2372
rect 4804 2320 4856 2372
rect 3792 2252 3844 2304
rect 7012 2252 7064 2304
rect 8300 2252 8352 2304
rect 9588 2252 9640 2304
rect 10600 2252 10652 2304
rect 12164 2252 12216 2304
rect 13452 2252 13504 2304
rect 14740 2252 14792 2304
rect 16028 2252 16080 2304
rect 17316 2252 17368 2304
rect 18880 2252 18932 2304
rect 5848 2150 5900 2202
rect 5912 2150 5964 2202
rect 5976 2150 6028 2202
rect 6040 2150 6092 2202
rect 6104 2150 6156 2202
rect 10747 2150 10799 2202
rect 10811 2150 10863 2202
rect 10875 2150 10927 2202
rect 10939 2150 10991 2202
rect 11003 2150 11055 2202
rect 15646 2150 15698 2202
rect 15710 2150 15762 2202
rect 15774 2150 15826 2202
rect 15838 2150 15890 2202
rect 15902 2150 15954 2202
rect 20545 2150 20597 2202
rect 20609 2150 20661 2202
rect 20673 2150 20725 2202
rect 20737 2150 20789 2202
rect 20801 2150 20853 2202
<< metal2 >>
rect 570 23205 626 24005
rect 1858 23205 1914 24005
rect 3146 23205 3202 24005
rect 4434 23338 4490 24005
rect 4434 23310 4660 23338
rect 4434 23205 4490 23310
rect 584 21146 612 23205
rect 1674 21856 1730 21865
rect 1674 21791 1730 21800
rect 572 21140 624 21146
rect 572 21082 624 21088
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1100 18540 1480 18560
rect 1100 18460 1120 18540
rect 1470 18460 1480 18540
rect 1100 18440 1480 18460
rect 1596 17338 1624 20878
rect 1688 20602 1716 21791
rect 1872 21690 1900 23205
rect 3160 21690 3188 23205
rect 4632 21690 4660 23310
rect 5722 23205 5778 24005
rect 7010 23338 7066 24005
rect 7010 23310 7328 23338
rect 7010 23205 7066 23310
rect 5736 21690 5764 23205
rect 5848 21788 6156 21797
rect 5848 21786 5854 21788
rect 5910 21786 5934 21788
rect 5990 21786 6014 21788
rect 6070 21786 6094 21788
rect 6150 21786 6156 21788
rect 5910 21734 5912 21786
rect 6092 21734 6094 21786
rect 5848 21732 5854 21734
rect 5910 21732 5934 21734
rect 5990 21732 6014 21734
rect 6070 21732 6094 21734
rect 6150 21732 6156 21734
rect 5848 21723 6156 21732
rect 7300 21690 7328 23310
rect 8298 23205 8354 24005
rect 9586 23205 9642 24005
rect 10874 23338 10930 24005
rect 10612 23310 10930 23338
rect 8312 21690 8340 23205
rect 9600 21706 9628 23205
rect 9600 21690 9720 21706
rect 10612 21690 10640 23310
rect 10874 23205 10930 23310
rect 12162 23338 12218 24005
rect 13450 23338 13506 24005
rect 12162 23310 12388 23338
rect 12162 23205 12218 23310
rect 10747 21788 11055 21797
rect 10747 21786 10753 21788
rect 10809 21786 10833 21788
rect 10889 21786 10913 21788
rect 10969 21786 10993 21788
rect 11049 21786 11055 21788
rect 10809 21734 10811 21786
rect 10991 21734 10993 21786
rect 10747 21732 10753 21734
rect 10809 21732 10833 21734
rect 10889 21732 10913 21734
rect 10969 21732 10993 21734
rect 11049 21732 11055 21734
rect 10747 21723 11055 21732
rect 12360 21690 12388 23310
rect 13450 23310 13768 23338
rect 13450 23205 13506 23310
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 8300 21684 8352 21690
rect 9600 21684 9732 21690
rect 9600 21678 9680 21684
rect 8300 21626 8352 21632
rect 9680 21626 9732 21632
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 12348 21684 12400 21690
rect 13740 21672 13768 23310
rect 14738 23205 14794 24005
rect 16026 23205 16082 24005
rect 17314 23205 17370 24005
rect 18602 23205 18658 24005
rect 19890 23205 19946 24005
rect 21178 23205 21234 24005
rect 14752 21690 14780 23205
rect 15646 21788 15954 21797
rect 15646 21786 15652 21788
rect 15708 21786 15732 21788
rect 15788 21786 15812 21788
rect 15868 21786 15892 21788
rect 15948 21786 15954 21788
rect 15708 21734 15710 21786
rect 15890 21734 15892 21786
rect 15646 21732 15652 21734
rect 15708 21732 15732 21734
rect 15788 21732 15812 21734
rect 15868 21732 15892 21734
rect 15948 21732 15954 21734
rect 15646 21723 15954 21732
rect 16040 21690 16068 23205
rect 16486 22672 16542 22681
rect 16486 22607 16542 22616
rect 13820 21684 13872 21690
rect 13740 21644 13820 21672
rect 12348 21626 12400 21632
rect 13820 21626 13872 21632
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2608 19446 2636 20402
rect 2700 20058 2728 20878
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2792 20534 2820 20810
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2792 19854 2820 20198
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2332 18834 2360 19246
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 18290 2360 18770
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17678 1992 18022
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 2516 16658 2544 17478
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15706 1992 15982
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1492 15496 1544 15502
rect 1492 15438 1544 15444
rect 1504 13938 1532 15438
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 13977 1624 14962
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 14414 1900 14758
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1582 13968 1638 13977
rect 1492 13932 1544 13938
rect 1582 13903 1638 13912
rect 1492 13874 1544 13880
rect 1504 13462 1532 13874
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12238 1624 12582
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1504 6914 1532 11222
rect 1780 11150 1808 12038
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10033 1624 10610
rect 1676 10056 1728 10062
rect 1582 10024 1638 10033
rect 1676 9998 1728 10004
rect 1582 9959 1638 9968
rect 1688 9518 1716 9998
rect 1872 9586 1900 14350
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1964 13326 1992 14214
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 2056 12850 2084 16594
rect 2608 16250 2636 17206
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1964 9518 1992 10406
rect 2332 10266 2360 10610
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2516 8634 2544 15982
rect 2700 15502 2728 17614
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3068 17270 3096 17478
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13326 2912 14214
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10062 2820 10406
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 7206 1716 7822
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6934 1716 7142
rect 1676 6928 1728 6934
rect 1504 6886 1624 6914
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 584 800 612 3606
rect 1596 3534 1624 6886
rect 1676 6870 1728 6876
rect 1872 6254 1900 7278
rect 2332 6798 2360 7686
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 2516 5370 2544 7414
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2516 4554 2544 5306
rect 2792 4690 2820 8570
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 6458 2912 8298
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2884 5710 2912 6258
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1688 3058 1716 4422
rect 2516 4214 2544 4490
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1780 2145 1808 3334
rect 2332 3058 2360 3878
rect 2516 3194 2544 4150
rect 2976 3942 3004 9454
rect 3160 9042 3188 17206
rect 3252 16250 3280 21490
rect 3399 21244 3707 21253
rect 3399 21242 3405 21244
rect 3461 21242 3485 21244
rect 3541 21242 3565 21244
rect 3621 21242 3645 21244
rect 3701 21242 3707 21244
rect 3461 21190 3463 21242
rect 3643 21190 3645 21242
rect 3399 21188 3405 21190
rect 3461 21188 3485 21190
rect 3541 21188 3565 21190
rect 3621 21188 3645 21190
rect 3701 21188 3707 21190
rect 3399 21179 3707 21188
rect 3884 20868 3936 20874
rect 3884 20810 3936 20816
rect 3399 20156 3707 20165
rect 3399 20154 3405 20156
rect 3461 20154 3485 20156
rect 3541 20154 3565 20156
rect 3621 20154 3645 20156
rect 3701 20154 3707 20156
rect 3461 20102 3463 20154
rect 3643 20102 3645 20154
rect 3399 20100 3405 20102
rect 3461 20100 3485 20102
rect 3541 20100 3565 20102
rect 3621 20100 3645 20102
rect 3701 20100 3707 20102
rect 3399 20091 3707 20100
rect 3399 19068 3707 19077
rect 3399 19066 3405 19068
rect 3461 19066 3485 19068
rect 3541 19066 3565 19068
rect 3621 19066 3645 19068
rect 3701 19066 3707 19068
rect 3461 19014 3463 19066
rect 3643 19014 3645 19066
rect 3399 19012 3405 19014
rect 3461 19012 3485 19014
rect 3541 19012 3565 19014
rect 3621 19012 3645 19014
rect 3701 19012 3707 19014
rect 3399 19003 3707 19012
rect 3399 17980 3707 17989
rect 3399 17978 3405 17980
rect 3461 17978 3485 17980
rect 3541 17978 3565 17980
rect 3621 17978 3645 17980
rect 3701 17978 3707 17980
rect 3461 17926 3463 17978
rect 3643 17926 3645 17978
rect 3399 17924 3405 17926
rect 3461 17924 3485 17926
rect 3541 17924 3565 17926
rect 3621 17924 3645 17926
rect 3701 17924 3707 17926
rect 3399 17915 3707 17924
rect 3896 17202 3924 20810
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3399 16892 3707 16901
rect 3399 16890 3405 16892
rect 3461 16890 3485 16892
rect 3541 16890 3565 16892
rect 3621 16890 3645 16892
rect 3701 16890 3707 16892
rect 3461 16838 3463 16890
rect 3643 16838 3645 16890
rect 3399 16836 3405 16838
rect 3461 16836 3485 16838
rect 3541 16836 3565 16838
rect 3621 16836 3645 16838
rect 3701 16836 3707 16838
rect 3399 16827 3707 16836
rect 3896 16590 3924 17138
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 16658 4016 16934
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3399 15804 3707 15813
rect 3399 15802 3405 15804
rect 3461 15802 3485 15804
rect 3541 15802 3565 15804
rect 3621 15802 3645 15804
rect 3701 15802 3707 15804
rect 3461 15750 3463 15802
rect 3643 15750 3645 15802
rect 3399 15748 3405 15750
rect 3461 15748 3485 15750
rect 3541 15748 3565 15750
rect 3621 15748 3645 15750
rect 3701 15748 3707 15750
rect 3399 15739 3707 15748
rect 3399 14716 3707 14725
rect 3399 14714 3405 14716
rect 3461 14714 3485 14716
rect 3541 14714 3565 14716
rect 3621 14714 3645 14716
rect 3701 14714 3707 14716
rect 3461 14662 3463 14714
rect 3643 14662 3645 14714
rect 3399 14660 3405 14662
rect 3461 14660 3485 14662
rect 3541 14660 3565 14662
rect 3621 14660 3645 14662
rect 3701 14660 3707 14662
rect 3399 14651 3707 14660
rect 3804 14006 3832 16118
rect 4080 14074 4108 21490
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4264 20262 4292 20470
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4264 19446 4292 20198
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 4264 19258 4292 19382
rect 4264 19230 4384 19258
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18834 4292 19110
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4356 18698 4384 19230
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 17746 4200 18022
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4540 17610 4568 18226
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 4540 16658 4568 17546
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4540 14074 4568 14282
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 3399 13628 3707 13637
rect 3399 13626 3405 13628
rect 3461 13626 3485 13628
rect 3541 13626 3565 13628
rect 3621 13626 3645 13628
rect 3701 13626 3707 13628
rect 3461 13574 3463 13626
rect 3643 13574 3645 13626
rect 3399 13572 3405 13574
rect 3461 13572 3485 13574
rect 3541 13572 3565 13574
rect 3621 13572 3645 13574
rect 3701 13572 3707 13574
rect 3399 13563 3707 13572
rect 4724 13530 4752 13874
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 3399 12540 3707 12549
rect 3399 12538 3405 12540
rect 3461 12538 3485 12540
rect 3541 12538 3565 12540
rect 3621 12538 3645 12540
rect 3701 12538 3707 12540
rect 3461 12486 3463 12538
rect 3643 12486 3645 12538
rect 3399 12484 3405 12486
rect 3461 12484 3485 12486
rect 3541 12484 3565 12486
rect 3621 12484 3645 12486
rect 3701 12484 3707 12486
rect 3399 12475 3707 12484
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11762 3556 12038
rect 4356 11898 4384 12786
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3399 11452 3707 11461
rect 3399 11450 3405 11452
rect 3461 11450 3485 11452
rect 3541 11450 3565 11452
rect 3621 11450 3645 11452
rect 3701 11450 3707 11452
rect 3461 11398 3463 11450
rect 3643 11398 3645 11450
rect 3399 11396 3405 11398
rect 3461 11396 3485 11398
rect 3541 11396 3565 11398
rect 3621 11396 3645 11398
rect 3701 11396 3707 11398
rect 3399 11387 3707 11396
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10810 4016 11086
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3252 10266 3280 10610
rect 3399 10364 3707 10373
rect 3399 10362 3405 10364
rect 3461 10362 3485 10364
rect 3541 10362 3565 10364
rect 3621 10362 3645 10364
rect 3701 10362 3707 10364
rect 3461 10310 3463 10362
rect 3643 10310 3645 10362
rect 3399 10308 3405 10310
rect 3461 10308 3485 10310
rect 3541 10308 3565 10310
rect 3621 10308 3645 10310
rect 3701 10308 3707 10310
rect 3399 10299 3707 10308
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 4540 9518 4568 13262
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11898 4844 12174
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4632 11354 4660 11698
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4908 9654 4936 21490
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 19922 5580 20742
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5644 19122 5672 21490
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 5848 20700 6156 20709
rect 5848 20698 5854 20700
rect 5910 20698 5934 20700
rect 5990 20698 6014 20700
rect 6070 20698 6094 20700
rect 6150 20698 6156 20700
rect 5910 20646 5912 20698
rect 6092 20646 6094 20698
rect 5848 20644 5854 20646
rect 5910 20644 5934 20646
rect 5990 20644 6014 20646
rect 6070 20644 6094 20646
rect 6150 20644 6156 20646
rect 5848 20635 6156 20644
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5736 19854 5764 20334
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 6564 19786 6592 20878
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6932 20618 6960 20810
rect 6932 20590 7052 20618
rect 7024 20262 7052 20590
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7024 19786 7052 20198
rect 7300 20058 7328 20402
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 5848 19612 6156 19621
rect 5848 19610 5854 19612
rect 5910 19610 5934 19612
rect 5990 19610 6014 19612
rect 6070 19610 6094 19612
rect 6150 19610 6156 19612
rect 5910 19558 5912 19610
rect 6092 19558 6094 19610
rect 5848 19556 5854 19558
rect 5910 19556 5934 19558
rect 5990 19556 6014 19558
rect 6070 19556 6094 19558
rect 6150 19556 6156 19558
rect 5848 19547 6156 19556
rect 5644 19094 5764 19122
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5092 18222 5120 18566
rect 5644 18358 5672 18566
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5092 17678 5120 18158
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5644 15094 5672 16390
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5368 14346 5396 14962
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 14074 5396 14282
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5552 13394 5580 14758
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12238 5212 12582
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5276 11150 5304 12038
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 3252 9178 3280 9454
rect 3399 9276 3707 9285
rect 3399 9274 3405 9276
rect 3461 9274 3485 9276
rect 3541 9274 3565 9276
rect 3621 9274 3645 9276
rect 3701 9274 3707 9276
rect 3461 9222 3463 9274
rect 3643 9222 3645 9274
rect 3399 9220 3405 9222
rect 3461 9220 3485 9222
rect 3541 9220 3565 9222
rect 3621 9220 3645 9222
rect 3701 9220 3707 9222
rect 3399 9211 3707 9220
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 4540 8974 4568 9454
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 3160 7886 3188 8366
rect 3399 8188 3707 8197
rect 3399 8186 3405 8188
rect 3461 8186 3485 8188
rect 3541 8186 3565 8188
rect 3621 8186 3645 8188
rect 3701 8186 3707 8188
rect 3461 8134 3463 8186
rect 3643 8134 3645 8186
rect 3399 8132 3405 8134
rect 3461 8132 3485 8134
rect 3541 8132 3565 8134
rect 3621 8132 3645 8134
rect 3701 8132 3707 8134
rect 3399 8123 3707 8132
rect 4264 8090 4292 8366
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7002 3188 7822
rect 3252 7206 3280 7958
rect 4356 7886 4384 8774
rect 5276 8634 5304 8842
rect 5264 8628 5316 8634
rect 5316 8588 5396 8616
rect 5264 8570 5316 8576
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3252 6322 3280 7142
rect 3399 7100 3707 7109
rect 3399 7098 3405 7100
rect 3461 7098 3485 7100
rect 3541 7098 3565 7100
rect 3621 7098 3645 7100
rect 3701 7098 3707 7100
rect 3461 7046 3463 7098
rect 3643 7046 3645 7098
rect 3399 7044 3405 7046
rect 3461 7044 3485 7046
rect 3541 7044 3565 7046
rect 3621 7044 3645 7046
rect 3701 7044 3707 7046
rect 3399 7035 3707 7044
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3804 6254 3832 7142
rect 3988 6798 4016 7686
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4356 7002 4384 7210
rect 4816 7206 4844 8502
rect 5368 8362 5396 8588
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3160 5778 3188 6190
rect 3399 6012 3707 6021
rect 3399 6010 3405 6012
rect 3461 6010 3485 6012
rect 3541 6010 3565 6012
rect 3621 6010 3645 6012
rect 3701 6010 3707 6012
rect 3461 5958 3463 6010
rect 3643 5958 3645 6010
rect 3399 5956 3405 5958
rect 3461 5956 3485 5958
rect 3541 5956 3565 5958
rect 3621 5956 3645 5958
rect 3701 5956 3707 5958
rect 3399 5947 3707 5956
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3160 4622 3188 5714
rect 3988 5710 4016 6258
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4540 5234 4568 6054
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5370 4752 5578
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 3399 4924 3707 4933
rect 3399 4922 3405 4924
rect 3461 4922 3485 4924
rect 3541 4922 3565 4924
rect 3621 4922 3645 4924
rect 3701 4922 3707 4924
rect 3461 4870 3463 4922
rect 3643 4870 3645 4922
rect 3399 4868 3405 4870
rect 3461 4868 3485 4870
rect 3541 4868 3565 4870
rect 3621 4868 3645 4870
rect 3701 4868 3707 4870
rect 3399 4859 3707 4868
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3160 4146 3188 4558
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1766 2136 1822 2145
rect 1766 2071 1822 2080
rect 1872 800 1900 2790
rect 2516 2378 2544 3130
rect 2976 3058 3004 3878
rect 3160 3058 3188 4082
rect 3399 3836 3707 3845
rect 3399 3834 3405 3836
rect 3461 3834 3485 3836
rect 3541 3834 3565 3836
rect 3621 3834 3645 3836
rect 3701 3834 3707 3836
rect 3461 3782 3463 3834
rect 3643 3782 3645 3834
rect 3399 3780 3405 3782
rect 3461 3780 3485 3782
rect 3541 3780 3565 3782
rect 3621 3780 3645 3782
rect 3701 3780 3707 3782
rect 3399 3771 3707 3780
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 3068 1442 3096 2790
rect 3252 2650 3280 3470
rect 4264 2990 4292 3538
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3399 2748 3707 2757
rect 3399 2746 3405 2748
rect 3461 2746 3485 2748
rect 3541 2746 3565 2748
rect 3621 2746 3645 2748
rect 3701 2746 3707 2748
rect 3461 2694 3463 2746
rect 3643 2694 3645 2746
rect 3399 2692 3405 2694
rect 3461 2692 3485 2694
rect 3541 2692 3565 2694
rect 3621 2692 3645 2694
rect 3701 2692 3707 2694
rect 3399 2683 3707 2692
rect 3804 2650 3832 2926
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3804 2310 3832 2586
rect 4264 2378 4292 2926
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3068 1414 3188 1442
rect 3160 800 3188 1414
rect 4448 800 4476 3334
rect 4632 3194 4660 3470
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4816 2378 4844 7142
rect 5368 6798 5396 8298
rect 5460 7954 5488 8842
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5552 7342 5580 9522
rect 5736 8634 5764 19094
rect 6564 18766 6592 19722
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 5848 18524 6156 18533
rect 5848 18522 5854 18524
rect 5910 18522 5934 18524
rect 5990 18522 6014 18524
rect 6070 18522 6094 18524
rect 6150 18522 6156 18524
rect 5910 18470 5912 18522
rect 6092 18470 6094 18522
rect 5848 18468 5854 18470
rect 5910 18468 5934 18470
rect 5990 18468 6014 18470
rect 6070 18468 6094 18470
rect 6150 18468 6156 18470
rect 5848 18459 6156 18468
rect 6564 18222 6592 18702
rect 7024 18630 7052 19722
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18426 7052 18566
rect 7116 18426 7144 18634
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17882 6868 18158
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 5848 17436 6156 17445
rect 5848 17434 5854 17436
rect 5910 17434 5934 17436
rect 5990 17434 6014 17436
rect 6070 17434 6094 17436
rect 6150 17434 6156 17436
rect 5910 17382 5912 17434
rect 6092 17382 6094 17434
rect 5848 17380 5854 17382
rect 5910 17380 5934 17382
rect 5990 17380 6014 17382
rect 6070 17380 6094 17382
rect 6150 17380 6156 17382
rect 5848 17371 6156 17380
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 16658 6868 16934
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 5848 16348 6156 16357
rect 5848 16346 5854 16348
rect 5910 16346 5934 16348
rect 5990 16346 6014 16348
rect 6070 16346 6094 16348
rect 6150 16346 6156 16348
rect 5910 16294 5912 16346
rect 6092 16294 6094 16346
rect 5848 16292 5854 16294
rect 5910 16292 5934 16294
rect 5990 16292 6014 16294
rect 6070 16292 6094 16294
rect 6150 16292 6156 16294
rect 5848 16283 6156 16292
rect 7300 16250 7328 17138
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6840 15502 6868 16050
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 5848 15260 6156 15269
rect 5848 15258 5854 15260
rect 5910 15258 5934 15260
rect 5990 15258 6014 15260
rect 6070 15258 6094 15260
rect 6150 15258 6156 15260
rect 5910 15206 5912 15258
rect 6092 15206 6094 15258
rect 5848 15204 5854 15206
rect 5910 15204 5934 15206
rect 5990 15204 6014 15206
rect 6070 15204 6094 15206
rect 6150 15204 6156 15206
rect 5848 15195 6156 15204
rect 5848 14172 6156 14181
rect 5848 14170 5854 14172
rect 5910 14170 5934 14172
rect 5990 14170 6014 14172
rect 6070 14170 6094 14172
rect 6150 14170 6156 14172
rect 5910 14118 5912 14170
rect 6092 14118 6094 14170
rect 5848 14116 5854 14118
rect 5910 14116 5934 14118
rect 5990 14116 6014 14118
rect 6070 14116 6094 14118
rect 6150 14116 6156 14118
rect 5848 14107 6156 14116
rect 6840 13938 6868 15438
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 14822 7328 15370
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14346 7328 14758
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13938 7236 14214
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 5848 13084 6156 13093
rect 5848 13082 5854 13084
rect 5910 13082 5934 13084
rect 5990 13082 6014 13084
rect 6070 13082 6094 13084
rect 6150 13082 6156 13084
rect 5910 13030 5912 13082
rect 6092 13030 6094 13082
rect 5848 13028 5854 13030
rect 5910 13028 5934 13030
rect 5990 13028 6014 13030
rect 6070 13028 6094 13030
rect 6150 13028 6156 13030
rect 5848 13019 6156 13028
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5848 11996 6156 12005
rect 5848 11994 5854 11996
rect 5910 11994 5934 11996
rect 5990 11994 6014 11996
rect 6070 11994 6094 11996
rect 6150 11994 6156 11996
rect 5910 11942 5912 11994
rect 6092 11942 6094 11994
rect 5848 11940 5854 11942
rect 5910 11940 5934 11942
rect 5990 11940 6014 11942
rect 6070 11940 6094 11942
rect 6150 11940 6156 11942
rect 5848 11931 6156 11940
rect 6196 11762 6224 12174
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11218 6224 11494
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 5848 10908 6156 10917
rect 5848 10906 5854 10908
rect 5910 10906 5934 10908
rect 5990 10906 6014 10908
rect 6070 10906 6094 10908
rect 6150 10906 6156 10908
rect 5910 10854 5912 10906
rect 6092 10854 6094 10906
rect 5848 10852 5854 10854
rect 5910 10852 5934 10854
rect 5990 10852 6014 10854
rect 6070 10852 6094 10854
rect 6150 10852 6156 10854
rect 5848 10843 6156 10852
rect 5848 9820 6156 9829
rect 5848 9818 5854 9820
rect 5910 9818 5934 9820
rect 5990 9818 6014 9820
rect 6070 9818 6094 9820
rect 6150 9818 6156 9820
rect 5910 9766 5912 9818
rect 6092 9766 6094 9818
rect 5848 9764 5854 9766
rect 5910 9764 5934 9766
rect 5990 9764 6014 9766
rect 6070 9764 6094 9766
rect 6150 9764 6156 9766
rect 5848 9755 6156 9764
rect 5848 8732 6156 8741
rect 5848 8730 5854 8732
rect 5910 8730 5934 8732
rect 5990 8730 6014 8732
rect 6070 8730 6094 8732
rect 6150 8730 6156 8732
rect 5910 8678 5912 8730
rect 6092 8678 6094 8730
rect 5848 8676 5854 8678
rect 5910 8676 5934 8678
rect 5990 8676 6014 8678
rect 6070 8676 6094 8678
rect 6150 8676 6156 8678
rect 5848 8667 6156 8676
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7410 5672 7822
rect 5848 7644 6156 7653
rect 5848 7642 5854 7644
rect 5910 7642 5934 7644
rect 5990 7642 6014 7644
rect 6070 7642 6094 7644
rect 6150 7642 6156 7644
rect 5910 7590 5912 7642
rect 6092 7590 6094 7642
rect 5848 7588 5854 7590
rect 5910 7588 5934 7590
rect 5990 7588 6014 7590
rect 6070 7588 6094 7590
rect 6150 7588 6156 7590
rect 5848 7579 6156 7588
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 6866 5672 7142
rect 5736 6866 5764 7278
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5356 6792 5408 6798
rect 5408 6752 5488 6780
rect 5356 6734 5408 6740
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5574 5120 6122
rect 5276 5846 5304 6190
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5092 4622 5120 5510
rect 5276 5370 5304 5782
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5460 4622 5488 6752
rect 5848 6556 6156 6565
rect 5848 6554 5854 6556
rect 5910 6554 5934 6556
rect 5990 6554 6014 6556
rect 6070 6554 6094 6556
rect 6150 6554 6156 6556
rect 5910 6502 5912 6554
rect 6092 6502 6094 6554
rect 5848 6500 5854 6502
rect 5910 6500 5934 6502
rect 5990 6500 6014 6502
rect 6070 6500 6094 6502
rect 6150 6500 6156 6502
rect 5848 6491 6156 6500
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5234 5672 6054
rect 6472 5914 6500 13806
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12442 6592 12718
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6840 12238 6868 13874
rect 7208 13394 7236 13874
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7300 13326 7328 14282
rect 7392 14074 7420 14350
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12918 7144 13126
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7116 12238 7144 12854
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6840 11898 6868 12174
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11354 6868 11698
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 9654 6868 11290
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8974 7328 9318
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7546 6868 7822
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5848 5468 6156 5477
rect 5848 5466 5854 5468
rect 5910 5466 5934 5468
rect 5990 5466 6014 5468
rect 6070 5466 6094 5468
rect 6150 5466 6156 5468
rect 5910 5414 5912 5466
rect 6092 5414 6094 5466
rect 5848 5412 5854 5414
rect 5910 5412 5934 5414
rect 5990 5412 6014 5414
rect 6070 5412 6094 5414
rect 6150 5412 6156 5414
rect 5848 5403 6156 5412
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 6196 4826 6224 5714
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 3602 5488 4558
rect 5848 4380 6156 4389
rect 5848 4378 5854 4380
rect 5910 4378 5934 4380
rect 5990 4378 6014 4380
rect 6070 4378 6094 4380
rect 6150 4378 6156 4380
rect 5910 4326 5912 4378
rect 6092 4326 6094 4378
rect 5848 4324 5854 4326
rect 5910 4324 5934 4326
rect 5990 4324 6014 4326
rect 6070 4324 6094 4326
rect 6150 4324 6156 4326
rect 5848 4315 6156 4324
rect 6472 4146 6500 5850
rect 6932 5370 6960 8842
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 7290 7328 7346
rect 7392 7290 7420 10542
rect 7484 9178 7512 21490
rect 8298 21244 8606 21253
rect 8298 21242 8304 21244
rect 8360 21242 8384 21244
rect 8440 21242 8464 21244
rect 8520 21242 8544 21244
rect 8600 21242 8606 21244
rect 8360 21190 8362 21242
rect 8542 21190 8544 21242
rect 8298 21188 8304 21190
rect 8360 21188 8384 21190
rect 8440 21188 8464 21190
rect 8520 21188 8544 21190
rect 8600 21188 8606 21190
rect 8298 21179 8606 21188
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8312 20466 8340 20742
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8036 19718 8064 20402
rect 8298 20156 8606 20165
rect 8298 20154 8304 20156
rect 8360 20154 8384 20156
rect 8440 20154 8464 20156
rect 8520 20154 8544 20156
rect 8600 20154 8606 20156
rect 8360 20102 8362 20154
rect 8542 20102 8544 20154
rect 8298 20100 8304 20102
rect 8360 20100 8384 20102
rect 8440 20100 8464 20102
rect 8520 20100 8544 20102
rect 8600 20100 8606 20102
rect 8298 20091 8606 20100
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 8036 19446 8064 19654
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8298 19068 8606 19077
rect 8298 19066 8304 19068
rect 8360 19066 8384 19068
rect 8440 19066 8464 19068
rect 8520 19066 8544 19068
rect 8600 19066 8606 19068
rect 8360 19014 8362 19066
rect 8542 19014 8544 19066
rect 8298 19012 8304 19014
rect 8360 19012 8384 19014
rect 8440 19012 8464 19014
rect 8520 19012 8544 19014
rect 8600 19012 8606 19014
rect 8298 19003 8606 19012
rect 8680 18970 8708 19110
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7576 18358 7604 18634
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 8298 17980 8606 17989
rect 8298 17978 8304 17980
rect 8360 17978 8384 17980
rect 8440 17978 8464 17980
rect 8520 17978 8544 17980
rect 8600 17978 8606 17980
rect 8360 17926 8362 17978
rect 8542 17926 8544 17978
rect 8298 17924 8304 17926
rect 8360 17924 8384 17926
rect 8440 17924 8464 17926
rect 8520 17924 8544 17926
rect 8600 17924 8606 17926
rect 8298 17915 8606 17924
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17202 7972 17478
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 16658 7788 16934
rect 8298 16892 8606 16901
rect 8298 16890 8304 16892
rect 8360 16890 8384 16892
rect 8440 16890 8464 16892
rect 8520 16890 8544 16892
rect 8600 16890 8606 16892
rect 8360 16838 8362 16890
rect 8542 16838 8544 16890
rect 8298 16836 8304 16838
rect 8360 16836 8384 16838
rect 8440 16836 8464 16838
rect 8520 16836 8544 16838
rect 8600 16836 8606 16838
rect 8298 16827 8606 16836
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8128 15434 8156 16458
rect 8680 16182 8708 16730
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8298 15804 8606 15813
rect 8298 15802 8304 15804
rect 8360 15802 8384 15804
rect 8440 15802 8464 15804
rect 8520 15802 8544 15804
rect 8600 15802 8606 15804
rect 8360 15750 8362 15802
rect 8542 15750 8544 15802
rect 8298 15748 8304 15750
rect 8360 15748 8384 15750
rect 8440 15748 8464 15750
rect 8520 15748 8544 15750
rect 8600 15748 8606 15750
rect 8298 15739 8606 15748
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7576 12918 7604 14826
rect 8128 13870 8156 15098
rect 8298 14716 8606 14725
rect 8298 14714 8304 14716
rect 8360 14714 8384 14716
rect 8440 14714 8464 14716
rect 8520 14714 8544 14716
rect 8600 14714 8606 14716
rect 8360 14662 8362 14714
rect 8542 14662 8544 14714
rect 8298 14660 8304 14662
rect 8360 14660 8384 14662
rect 8440 14660 8464 14662
rect 8520 14660 8544 14662
rect 8600 14660 8606 14662
rect 8298 14651 8606 14660
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8498 7512 8774
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7484 7410 7512 8434
rect 7576 8090 7604 12854
rect 7760 11082 7788 13194
rect 8128 12306 8156 13806
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8220 12238 8248 13874
rect 8772 13870 8800 14282
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8298 13628 8606 13637
rect 8298 13626 8304 13628
rect 8360 13626 8384 13628
rect 8440 13626 8464 13628
rect 8520 13626 8544 13628
rect 8600 13626 8606 13628
rect 8360 13574 8362 13626
rect 8542 13574 8544 13626
rect 8298 13572 8304 13574
rect 8360 13572 8384 13574
rect 8440 13572 8464 13574
rect 8520 13572 8544 13574
rect 8600 13572 8606 13574
rect 8298 13563 8606 13572
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8298 12540 8606 12549
rect 8298 12538 8304 12540
rect 8360 12538 8384 12540
rect 8440 12538 8464 12540
rect 8520 12538 8544 12540
rect 8600 12538 8606 12540
rect 8360 12486 8362 12538
rect 8542 12486 8544 12538
rect 8298 12484 8304 12486
rect 8360 12484 8384 12486
rect 8440 12484 8464 12486
rect 8520 12484 8544 12486
rect 8600 12484 8606 12486
rect 8298 12475 8606 12484
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11626 8248 12174
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 8128 8974 8156 11154
rect 8220 10674 8248 11562
rect 8298 11452 8606 11461
rect 8298 11450 8304 11452
rect 8360 11450 8384 11452
rect 8440 11450 8464 11452
rect 8520 11450 8544 11452
rect 8600 11450 8606 11452
rect 8360 11398 8362 11450
rect 8542 11398 8544 11450
rect 8298 11396 8304 11398
rect 8360 11396 8384 11398
rect 8440 11396 8464 11398
rect 8520 11396 8544 11398
rect 8600 11396 8606 11398
rect 8298 11387 8606 11396
rect 8680 11150 8708 12582
rect 8772 12442 8800 12786
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8298 10364 8606 10373
rect 8298 10362 8304 10364
rect 8360 10362 8384 10364
rect 8440 10362 8464 10364
rect 8520 10362 8544 10364
rect 8600 10362 8606 10364
rect 8360 10310 8362 10362
rect 8542 10310 8544 10362
rect 8298 10308 8304 10310
rect 8360 10308 8384 10310
rect 8440 10308 8464 10310
rect 8520 10308 8544 10310
rect 8600 10308 8606 10310
rect 8298 10299 8606 10308
rect 8680 10062 8708 10950
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8772 9926 8800 10678
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8298 9276 8606 9285
rect 8298 9274 8304 9276
rect 8360 9274 8384 9276
rect 8440 9274 8464 9276
rect 8520 9274 8544 9276
rect 8600 9274 8606 9276
rect 8360 9222 8362 9274
rect 8542 9222 8544 9274
rect 8298 9220 8304 9222
rect 8360 9220 8384 9222
rect 8440 9220 8464 9222
rect 8520 9220 8544 9222
rect 8600 9220 8606 9222
rect 8298 9211 8606 9220
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8566 7972 8774
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 8128 7954 8156 8910
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8298 8188 8606 8197
rect 8298 8186 8304 8188
rect 8360 8186 8384 8188
rect 8440 8186 8464 8188
rect 8520 8186 8544 8188
rect 8600 8186 8606 8188
rect 8360 8134 8362 8186
rect 8542 8134 8544 8186
rect 8298 8132 8304 8134
rect 8360 8132 8384 8134
rect 8440 8132 8464 8134
rect 8520 8132 8544 8134
rect 8600 8132 8606 8134
rect 8298 8123 8606 8132
rect 8680 8090 8708 8502
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8680 7410 8708 8026
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 7300 7262 7420 7290
rect 7392 6254 7420 7262
rect 8298 7100 8606 7109
rect 8298 7098 8304 7100
rect 8360 7098 8384 7100
rect 8440 7098 8464 7100
rect 8520 7098 8544 7100
rect 8600 7098 8606 7100
rect 8360 7046 8362 7098
rect 8542 7046 8544 7098
rect 8298 7044 8304 7046
rect 8360 7044 8384 7046
rect 8440 7044 8464 7046
rect 8520 7044 8544 7046
rect 8600 7044 8606 7046
rect 8298 7035 8606 7044
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7484 6458 7512 6666
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7484 6322 7512 6394
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6656 4282 6684 4490
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 6932 3466 6960 5306
rect 7392 4078 7420 6190
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5302 7880 6054
rect 7944 5846 7972 6598
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8298 6012 8606 6021
rect 8298 6010 8304 6012
rect 8360 6010 8384 6012
rect 8440 6010 8464 6012
rect 8520 6010 8544 6012
rect 8600 6010 8606 6012
rect 8360 5958 8362 6010
rect 8542 5958 8544 6010
rect 8298 5956 8304 5958
rect 8360 5956 8384 5958
rect 8440 5956 8464 5958
rect 8520 5956 8544 5958
rect 8600 5956 8606 5958
rect 8298 5947 8606 5956
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7944 5710 7972 5782
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7944 5166 7972 5646
rect 8772 5370 8800 6054
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8298 4924 8606 4933
rect 8298 4922 8304 4924
rect 8360 4922 8384 4924
rect 8440 4922 8464 4924
rect 8520 4922 8544 4924
rect 8600 4922 8606 4924
rect 8360 4870 8362 4922
rect 8542 4870 8544 4922
rect 8298 4868 8304 4870
rect 8360 4868 8384 4870
rect 8440 4868 8464 4870
rect 8520 4868 8544 4870
rect 8600 4868 8606 4870
rect 8298 4859 8606 4868
rect 8772 4690 8800 5306
rect 8956 4826 8984 21490
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9232 19378 9260 19858
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9508 17678 9536 20878
rect 9692 20602 9720 21490
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9864 20528 9916 20534
rect 9864 20470 9916 20476
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 17882 9720 18158
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17672 9548 17678
rect 9548 17620 9628 17626
rect 9496 17614 9628 17620
rect 9508 17598 9628 17614
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9508 16794 9536 17138
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9600 15162 9628 17598
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9692 17338 9720 17546
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9784 16114 9812 16458
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9784 15434 9812 16050
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9140 14482 9168 14894
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9876 14346 9904 20470
rect 10152 20466 10180 20878
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 16250 10088 16526
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9876 14006 9904 14282
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 12306 9168 12582
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9876 12170 9904 13942
rect 9968 13938 9996 14758
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9968 12646 9996 12786
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12306 9996 12582
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 10244 11082 10272 18158
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 6798 9168 7142
rect 9232 6866 9260 10542
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9586 9352 9862
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9508 8498 9536 11018
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10062 9628 10406
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9508 7818 9536 8434
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 7546 9536 7754
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9232 6322 9260 6802
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9416 5370 9444 5578
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 5166 9444 5306
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 5368 3126 5396 3402
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 5848 3292 6156 3301
rect 5848 3290 5854 3292
rect 5910 3290 5934 3292
rect 5990 3290 6014 3292
rect 6070 3290 6094 3292
rect 6150 3290 6156 3292
rect 5910 3238 5912 3290
rect 6092 3238 6094 3290
rect 5848 3236 5854 3238
rect 5910 3236 5934 3238
rect 5990 3236 6014 3238
rect 6070 3236 6094 3238
rect 6150 3236 6156 3238
rect 5848 3227 6156 3236
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5368 2650 5396 3062
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 5736 800 5764 2790
rect 6012 2650 6040 2994
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 7116 2446 7144 3334
rect 7944 3058 7972 4490
rect 8772 4214 8800 4626
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8220 2990 8248 4014
rect 8298 3836 8606 3845
rect 8298 3834 8304 3836
rect 8360 3834 8384 3836
rect 8440 3834 8464 3836
rect 8520 3834 8544 3836
rect 8600 3834 8606 3836
rect 8360 3782 8362 3834
rect 8542 3782 8544 3834
rect 8298 3780 8304 3782
rect 8360 3780 8384 3782
rect 8440 3780 8464 3782
rect 8520 3780 8544 3782
rect 8600 3780 8606 3782
rect 8298 3771 8606 3780
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8298 2748 8606 2757
rect 8298 2746 8304 2748
rect 8360 2746 8384 2748
rect 8440 2746 8464 2748
rect 8520 2746 8544 2748
rect 8600 2746 8606 2748
rect 8360 2694 8362 2746
rect 8542 2694 8544 2746
rect 8298 2692 8304 2694
rect 8360 2692 8384 2694
rect 8440 2692 8464 2694
rect 8520 2692 8544 2694
rect 8600 2692 8606 2694
rect 8298 2683 8606 2692
rect 8680 2446 8708 2790
rect 9600 2774 9628 8978
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9692 7478 9720 8230
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9692 6798 9720 7414
rect 9784 7342 9812 8774
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 3942 9720 6054
rect 9784 5778 9812 6122
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9772 3052 9824 3058
rect 9876 3040 9904 11018
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9968 9722 9996 9998
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10336 9466 10364 20334
rect 10428 19514 10456 20810
rect 10747 20700 11055 20709
rect 10747 20698 10753 20700
rect 10809 20698 10833 20700
rect 10889 20698 10913 20700
rect 10969 20698 10993 20700
rect 11049 20698 11055 20700
rect 10809 20646 10811 20698
rect 10991 20646 10993 20698
rect 10747 20644 10753 20646
rect 10809 20644 10833 20646
rect 10889 20644 10913 20646
rect 10969 20644 10993 20646
rect 11049 20644 11055 20646
rect 10747 20635 11055 20644
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11072 19922 11100 20402
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10747 19612 11055 19621
rect 10747 19610 10753 19612
rect 10809 19610 10833 19612
rect 10889 19610 10913 19612
rect 10969 19610 10993 19612
rect 11049 19610 11055 19612
rect 10809 19558 10811 19610
rect 10991 19558 10993 19610
rect 10747 19556 10753 19558
rect 10809 19556 10833 19558
rect 10889 19556 10913 19558
rect 10969 19556 10993 19558
rect 11049 19556 11055 19558
rect 10747 19547 11055 19556
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10747 18524 11055 18533
rect 10747 18522 10753 18524
rect 10809 18522 10833 18524
rect 10889 18522 10913 18524
rect 10969 18522 10993 18524
rect 11049 18522 11055 18524
rect 10809 18470 10811 18522
rect 10991 18470 10993 18522
rect 10747 18468 10753 18470
rect 10809 18468 10833 18470
rect 10889 18468 10913 18470
rect 10969 18468 10993 18470
rect 11049 18468 11055 18470
rect 10747 18459 11055 18468
rect 11164 18426 11192 21490
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11348 19922 11376 20742
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19530 11284 19654
rect 11440 19530 11468 20810
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 19854 12480 20198
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 11256 19502 11468 19530
rect 11256 19446 11284 19502
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11256 17882 11284 19382
rect 12544 18970 12572 21490
rect 13197 21244 13505 21253
rect 13197 21242 13203 21244
rect 13259 21242 13283 21244
rect 13339 21242 13363 21244
rect 13419 21242 13443 21244
rect 13499 21242 13505 21244
rect 13259 21190 13261 21242
rect 13441 21190 13443 21242
rect 13197 21188 13203 21190
rect 13259 21188 13283 21190
rect 13339 21188 13363 21190
rect 13419 21188 13443 21190
rect 13499 21188 13505 21190
rect 13197 21179 13505 21188
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13464 20602 13492 20878
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13464 20398 13492 20538
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 12820 20058 12848 20334
rect 13197 20156 13505 20165
rect 13197 20154 13203 20156
rect 13259 20154 13283 20156
rect 13339 20154 13363 20156
rect 13419 20154 13443 20156
rect 13499 20154 13505 20156
rect 13259 20102 13261 20154
rect 13441 20102 13443 20154
rect 13197 20100 13203 20102
rect 13259 20100 13283 20102
rect 13339 20100 13363 20102
rect 13419 20100 13443 20102
rect 13499 20100 13505 20102
rect 13197 20091 13505 20100
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 13197 19068 13505 19077
rect 13197 19066 13203 19068
rect 13259 19066 13283 19068
rect 13339 19066 13363 19068
rect 13419 19066 13443 19068
rect 13499 19066 13505 19068
rect 13259 19014 13261 19066
rect 13441 19014 13443 19066
rect 13197 19012 13203 19014
rect 13259 19012 13283 19014
rect 13339 19012 13363 19014
rect 13419 19012 13443 19014
rect 13499 19012 13505 19014
rect 13197 19003 13505 19012
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 10747 17436 11055 17445
rect 10747 17434 10753 17436
rect 10809 17434 10833 17436
rect 10889 17434 10913 17436
rect 10969 17434 10993 17436
rect 11049 17434 11055 17436
rect 10809 17382 10811 17434
rect 10991 17382 10993 17434
rect 10747 17380 10753 17382
rect 10809 17380 10833 17382
rect 10889 17380 10913 17382
rect 10969 17380 10993 17382
rect 11049 17380 11055 17382
rect 10747 17371 11055 17380
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 16046 10456 16594
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 10747 16348 11055 16357
rect 10747 16346 10753 16348
rect 10809 16346 10833 16348
rect 10889 16346 10913 16348
rect 10969 16346 10993 16348
rect 11049 16346 11055 16348
rect 10809 16294 10811 16346
rect 10991 16294 10993 16346
rect 10747 16292 10753 16294
rect 10809 16292 10833 16294
rect 10889 16292 10913 16294
rect 10969 16292 10993 16294
rect 11049 16292 11055 16294
rect 10747 16283 11055 16292
rect 11624 16114 11652 16390
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10520 15502 10548 16050
rect 11624 15570 11652 16050
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10747 15260 11055 15269
rect 10747 15258 10753 15260
rect 10809 15258 10833 15260
rect 10889 15258 10913 15260
rect 10969 15258 10993 15260
rect 11049 15258 11055 15260
rect 10809 15206 10811 15258
rect 10991 15206 10993 15258
rect 10747 15204 10753 15206
rect 10809 15204 10833 15206
rect 10889 15204 10913 15206
rect 10969 15204 10993 15206
rect 11049 15204 11055 15206
rect 10747 15195 11055 15204
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10888 14618 10916 14962
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10428 14074 10456 14418
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10428 13394 10456 14010
rect 10612 13462 10640 14554
rect 11164 14550 11192 14962
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14550 11376 14758
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11716 14278 11744 18566
rect 12084 18358 12112 18634
rect 12452 18426 12480 18770
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12452 18086 12480 18226
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17746 12480 18022
rect 13197 17980 13505 17989
rect 13197 17978 13203 17980
rect 13259 17978 13283 17980
rect 13339 17978 13363 17980
rect 13419 17978 13443 17980
rect 13499 17978 13505 17980
rect 13259 17926 13261 17978
rect 13441 17926 13443 17978
rect 13197 17924 13203 17926
rect 13259 17924 13283 17926
rect 13339 17924 13363 17926
rect 13419 17924 13443 17926
rect 13499 17924 13505 17926
rect 13197 17915 13505 17924
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 12452 16658 12480 17682
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12544 16794 12572 17138
rect 13197 16892 13505 16901
rect 13197 16890 13203 16892
rect 13259 16890 13283 16892
rect 13339 16890 13363 16892
rect 13419 16890 13443 16892
rect 13499 16890 13505 16892
rect 13259 16838 13261 16890
rect 13441 16838 13443 16890
rect 13197 16836 13203 16838
rect 13259 16836 13283 16838
rect 13339 16836 13363 16838
rect 13419 16836 13443 16838
rect 13499 16836 13505 16838
rect 13197 16827 13505 16836
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 13740 16522 13768 17614
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13197 15804 13505 15813
rect 13197 15802 13203 15804
rect 13259 15802 13283 15804
rect 13339 15802 13363 15804
rect 13419 15802 13443 15804
rect 13499 15802 13505 15804
rect 13259 15750 13261 15802
rect 13441 15750 13443 15802
rect 13197 15748 13203 15750
rect 13259 15748 13283 15750
rect 13339 15748 13363 15750
rect 13419 15748 13443 15750
rect 13499 15748 13505 15750
rect 13197 15739 13505 15748
rect 13740 15638 13768 16458
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 14108 15434 14136 17682
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12360 15026 12388 15302
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 14414 12296 14758
rect 12912 14414 12940 15098
rect 14108 15026 14136 15370
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 13197 14716 13505 14725
rect 13197 14714 13203 14716
rect 13259 14714 13283 14716
rect 13339 14714 13363 14716
rect 13419 14714 13443 14716
rect 13499 14714 13505 14716
rect 13259 14662 13261 14714
rect 13441 14662 13443 14714
rect 13197 14660 13203 14662
rect 13259 14660 13283 14662
rect 13339 14660 13363 14662
rect 13419 14660 13443 14662
rect 13499 14660 13505 14662
rect 13197 14651 13505 14660
rect 14108 14618 14136 14962
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 10747 14172 11055 14181
rect 10747 14170 10753 14172
rect 10809 14170 10833 14172
rect 10889 14170 10913 14172
rect 10969 14170 10993 14172
rect 11049 14170 11055 14172
rect 10809 14118 10811 14170
rect 10991 14118 10993 14170
rect 10747 14116 10753 14118
rect 10809 14116 10833 14118
rect 10889 14116 10913 14118
rect 10969 14116 10993 14118
rect 11049 14116 11055 14118
rect 10747 14107 11055 14116
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11072 13530 11100 13874
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10747 13084 11055 13093
rect 10747 13082 10753 13084
rect 10809 13082 10833 13084
rect 10889 13082 10913 13084
rect 10969 13082 10993 13084
rect 11049 13082 11055 13084
rect 10809 13030 10811 13082
rect 10991 13030 10993 13082
rect 10747 13028 10753 13030
rect 10809 13028 10833 13030
rect 10889 13028 10913 13030
rect 10969 13028 10993 13030
rect 11049 13028 11055 13030
rect 10747 13019 11055 13028
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10520 11762 10548 12582
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10747 11996 11055 12005
rect 10747 11994 10753 11996
rect 10809 11994 10833 11996
rect 10889 11994 10913 11996
rect 10969 11994 10993 11996
rect 11049 11994 11055 11996
rect 10809 11942 10811 11994
rect 10991 11942 10993 11994
rect 10747 11940 10753 11942
rect 10809 11940 10833 11942
rect 10889 11940 10913 11942
rect 10969 11940 10993 11942
rect 11049 11940 11055 11942
rect 10747 11931 11055 11940
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 11164 11694 11192 12378
rect 11256 11898 11284 12718
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 11286 10456 11494
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 11256 11218 11284 11834
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 10747 10908 11055 10917
rect 10747 10906 10753 10908
rect 10809 10906 10833 10908
rect 10889 10906 10913 10908
rect 10969 10906 10993 10908
rect 11049 10906 11055 10908
rect 10809 10854 10811 10906
rect 10991 10854 10993 10906
rect 10747 10852 10753 10854
rect 10809 10852 10833 10854
rect 10889 10852 10913 10854
rect 10969 10852 10993 10854
rect 11049 10852 11055 10854
rect 10747 10843 11055 10852
rect 11440 10266 11468 11086
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10520 9654 10548 9862
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10612 9586 10640 9998
rect 10747 9820 11055 9829
rect 10747 9818 10753 9820
rect 10809 9818 10833 9820
rect 10889 9818 10913 9820
rect 10969 9818 10993 9820
rect 11049 9818 11055 9820
rect 10809 9766 10811 9818
rect 10991 9766 10993 9818
rect 10747 9764 10753 9766
rect 10809 9764 10833 9766
rect 10889 9764 10913 9766
rect 10969 9764 10993 9766
rect 11049 9764 11055 9766
rect 10747 9755 11055 9764
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10336 9438 10456 9466
rect 10428 9382 10456 9438
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9968 8022 9996 8842
rect 10336 8498 10364 8910
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10336 8090 10364 8434
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 5914 9996 6190
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9968 5234 9996 5850
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10244 4622 10272 4966
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10428 4078 10456 9318
rect 10747 8732 11055 8741
rect 10747 8730 10753 8732
rect 10809 8730 10833 8732
rect 10889 8730 10913 8732
rect 10969 8730 10993 8732
rect 11049 8730 11055 8732
rect 10809 8678 10811 8730
rect 10991 8678 10993 8730
rect 10747 8676 10753 8678
rect 10809 8676 10833 8678
rect 10889 8676 10913 8678
rect 10969 8676 10993 8678
rect 11049 8676 11055 8678
rect 10747 8667 11055 8676
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10520 7954 10548 8230
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10747 7644 11055 7653
rect 10747 7642 10753 7644
rect 10809 7642 10833 7644
rect 10889 7642 10913 7644
rect 10969 7642 10993 7644
rect 11049 7642 11055 7644
rect 10809 7590 10811 7642
rect 10991 7590 10993 7642
rect 10747 7588 10753 7590
rect 10809 7588 10833 7590
rect 10889 7588 10913 7590
rect 10969 7588 10993 7590
rect 11049 7588 11055 7590
rect 10747 7579 11055 7588
rect 11164 7546 11192 8026
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6798 11468 7142
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10520 6118 10548 6326
rect 10612 6322 10640 6598
rect 10747 6556 11055 6565
rect 10747 6554 10753 6556
rect 10809 6554 10833 6556
rect 10889 6554 10913 6556
rect 10969 6554 10993 6556
rect 11049 6554 11055 6556
rect 10809 6502 10811 6554
rect 10991 6502 10993 6554
rect 10747 6500 10753 6502
rect 10809 6500 10833 6502
rect 10889 6500 10913 6502
rect 10969 6500 10993 6502
rect 11049 6500 11055 6502
rect 10747 6491 11055 6500
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5234 10548 6054
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10612 5166 10640 5578
rect 10747 5468 11055 5477
rect 10747 5466 10753 5468
rect 10809 5466 10833 5468
rect 10889 5466 10913 5468
rect 10969 5466 10993 5468
rect 11049 5466 11055 5468
rect 10809 5414 10811 5466
rect 10991 5414 10993 5466
rect 10747 5412 10753 5414
rect 10809 5412 10833 5414
rect 10889 5412 10913 5414
rect 10969 5412 10993 5414
rect 11049 5412 11055 5414
rect 10747 5403 11055 5412
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9824 3012 9904 3040
rect 9772 2994 9824 3000
rect 9508 2746 9628 2774
rect 9508 2514 9536 2746
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9968 2446 9996 3878
rect 10612 3670 10640 5102
rect 10747 4380 11055 4389
rect 10747 4378 10753 4380
rect 10809 4378 10833 4380
rect 10889 4378 10913 4380
rect 10969 4378 10993 4380
rect 11049 4378 11055 4380
rect 10809 4326 10811 4378
rect 10991 4326 10993 4378
rect 10747 4324 10753 4326
rect 10809 4324 10833 4326
rect 10889 4324 10913 4326
rect 10969 4324 10993 4326
rect 11049 4324 11055 4326
rect 10747 4315 11055 4324
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 11532 3602 11560 14214
rect 12544 13938 12572 14282
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12452 13462 12480 13806
rect 12820 13530 12848 13806
rect 13197 13628 13505 13637
rect 13197 13626 13203 13628
rect 13259 13626 13283 13628
rect 13339 13626 13363 13628
rect 13419 13626 13443 13628
rect 13499 13626 13505 13628
rect 13259 13574 13261 13626
rect 13441 13574 13443 13626
rect 13197 13572 13203 13574
rect 13259 13572 13283 13574
rect 13339 13572 13363 13574
rect 13419 13572 13443 13574
rect 13499 13572 13505 13574
rect 13197 13563 13505 13572
rect 14108 13530 14136 14554
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 13464 13326 13492 13466
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 12636 12782 12664 13262
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11716 12442 11744 12650
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 13096 12374 13124 13262
rect 13197 12540 13505 12549
rect 13197 12538 13203 12540
rect 13259 12538 13283 12540
rect 13339 12538 13363 12540
rect 13419 12538 13443 12540
rect 13499 12538 13505 12540
rect 13259 12486 13261 12538
rect 13441 12486 13443 12538
rect 13197 12484 13203 12486
rect 13259 12484 13283 12486
rect 13339 12484 13363 12486
rect 13419 12484 13443 12486
rect 13499 12484 13505 12486
rect 13197 12475 13505 12484
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11694 11744 12174
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 11992 11898 12020 12106
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10130 11652 10610
rect 11716 10606 11744 11630
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11900 10198 11928 10950
rect 12636 10742 12664 12106
rect 13096 11762 13124 12310
rect 13924 11830 13952 13262
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13197 11452 13505 11461
rect 13197 11450 13203 11452
rect 13259 11450 13283 11452
rect 13339 11450 13363 11452
rect 13419 11450 13443 11452
rect 13499 11450 13505 11452
rect 13259 11398 13261 11450
rect 13441 11398 13443 11450
rect 13197 11396 13203 11398
rect 13259 11396 13283 11398
rect 13339 11396 13363 11398
rect 13419 11396 13443 11398
rect 13499 11396 13505 11398
rect 13197 11387 13505 11396
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11992 9926 12020 10542
rect 12636 10266 12664 10678
rect 13924 10674 13952 11766
rect 14016 11694 14044 12106
rect 14108 12102 14136 12854
rect 14200 12442 14228 21490
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14292 20058 14320 21082
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14292 17746 14320 18158
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16114 14320 16526
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 13326 14320 14350
rect 14384 14074 14412 21490
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15764 21010 15792 21286
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 17882 14780 18158
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14660 16250 14688 17138
rect 15304 16250 15332 20878
rect 15646 20700 15954 20709
rect 15646 20698 15652 20700
rect 15708 20698 15732 20700
rect 15788 20698 15812 20700
rect 15868 20698 15892 20700
rect 15948 20698 15954 20700
rect 15708 20646 15710 20698
rect 15890 20646 15892 20698
rect 15646 20644 15652 20646
rect 15708 20644 15732 20646
rect 15788 20644 15812 20646
rect 15868 20644 15892 20646
rect 15948 20644 15954 20646
rect 15646 20635 15954 20644
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15396 20346 15424 20402
rect 16028 20392 16080 20398
rect 15396 20318 15516 20346
rect 16028 20334 16080 20340
rect 15488 20262 15516 20318
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15488 19786 15516 20198
rect 15764 19922 15792 20198
rect 16040 19922 16068 20334
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16500 19854 16528 22607
rect 17328 21690 17356 23205
rect 18616 21690 18644 23205
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15646 19612 15954 19621
rect 15646 19610 15652 19612
rect 15708 19610 15732 19612
rect 15788 19610 15812 19612
rect 15868 19610 15892 19612
rect 15948 19610 15954 19612
rect 15708 19558 15710 19610
rect 15890 19558 15892 19610
rect 15646 19556 15652 19558
rect 15708 19556 15732 19558
rect 15788 19556 15812 19558
rect 15868 19556 15892 19558
rect 15948 19556 15954 19558
rect 15646 19547 15954 19556
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16224 18834 16252 19314
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15396 18426 15424 18702
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15646 18524 15954 18533
rect 15646 18522 15652 18524
rect 15708 18522 15732 18524
rect 15788 18522 15812 18524
rect 15868 18522 15892 18524
rect 15948 18522 15954 18524
rect 15708 18470 15710 18522
rect 15890 18470 15892 18522
rect 15646 18468 15652 18470
rect 15708 18468 15732 18470
rect 15788 18468 15812 18470
rect 15868 18468 15892 18470
rect 15948 18468 15954 18470
rect 15646 18459 15954 18468
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15396 17338 15424 18362
rect 16040 18358 16068 18634
rect 16224 18426 16252 18770
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 15646 17436 15954 17445
rect 15646 17434 15652 17436
rect 15708 17434 15732 17436
rect 15788 17434 15812 17436
rect 15868 17434 15892 17436
rect 15948 17434 15954 17436
rect 15708 17382 15710 17434
rect 15890 17382 15892 17434
rect 15646 17380 15652 17382
rect 15708 17380 15732 17382
rect 15788 17380 15812 17382
rect 15868 17380 15892 17382
rect 15948 17380 15954 17382
rect 15646 17371 15954 17380
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 16040 17218 16068 18294
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 15948 17190 16068 17218
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15120 15570 15148 16050
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15304 15194 15332 16186
rect 15488 16114 15516 17070
rect 15948 16522 15976 17190
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 16040 16794 16068 17002
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15646 16348 15954 16357
rect 15646 16346 15652 16348
rect 15708 16346 15732 16348
rect 15788 16346 15812 16348
rect 15868 16346 15892 16348
rect 15948 16346 15954 16348
rect 15708 16294 15710 16346
rect 15890 16294 15892 16346
rect 15646 16292 15652 16294
rect 15708 16292 15732 16294
rect 15788 16292 15812 16294
rect 15868 16292 15892 16294
rect 15948 16292 15954 16294
rect 15646 16283 15954 16292
rect 16040 16114 16068 16730
rect 16500 16658 16528 17274
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16132 15434 16160 16458
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 15646 15260 15954 15269
rect 15646 15258 15652 15260
rect 15708 15258 15732 15260
rect 15788 15258 15812 15260
rect 15868 15258 15892 15260
rect 15948 15258 15954 15260
rect 15708 15206 15710 15258
rect 15890 15206 15892 15258
rect 15646 15204 15652 15206
rect 15708 15204 15732 15206
rect 15788 15204 15812 15206
rect 15868 15204 15892 15206
rect 15948 15204 15954 15206
rect 15646 15195 15954 15204
rect 15304 15166 15516 15194
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14482 14596 14758
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14660 12986 14688 13942
rect 15212 13394 15240 14282
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15212 13258 15240 13330
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14016 10588 14044 11630
rect 14188 10600 14240 10606
rect 14016 10560 14188 10588
rect 14188 10542 14240 10548
rect 13197 10364 13505 10373
rect 13197 10362 13203 10364
rect 13259 10362 13283 10364
rect 13339 10362 13363 10364
rect 13419 10362 13443 10364
rect 13499 10362 13505 10364
rect 13259 10310 13261 10362
rect 13441 10310 13443 10362
rect 13197 10308 13203 10310
rect 13259 10308 13283 10310
rect 13339 10308 13363 10310
rect 13419 10308 13443 10310
rect 13499 10308 13505 10310
rect 13197 10299 13505 10308
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9518 12020 9862
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 13197 9276 13505 9285
rect 13197 9274 13203 9276
rect 13259 9274 13283 9276
rect 13339 9274 13363 9276
rect 13419 9274 13443 9276
rect 13499 9274 13505 9276
rect 13259 9222 13261 9274
rect 13441 9222 13443 9274
rect 13197 9220 13203 9222
rect 13259 9220 13283 9222
rect 13339 9220 13363 9222
rect 13419 9220 13443 9222
rect 13499 9220 13505 9222
rect 13197 9211 13505 9220
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12084 8634 12112 8910
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12268 6934 12296 8978
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8566 12848 8774
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12912 7886 12940 8366
rect 13197 8188 13505 8197
rect 13197 8186 13203 8188
rect 13259 8186 13283 8188
rect 13339 8186 13363 8188
rect 13419 8186 13443 8188
rect 13499 8186 13505 8188
rect 13259 8134 13261 8186
rect 13441 8134 13443 8186
rect 13197 8132 13203 8134
rect 13259 8132 13283 8134
rect 13339 8132 13363 8134
rect 13419 8132 13443 8134
rect 13499 8132 13505 8134
rect 13197 8123 13505 8132
rect 13556 8090 13584 8910
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13556 7886 13584 8026
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13197 7100 13505 7109
rect 13197 7098 13203 7100
rect 13259 7098 13283 7100
rect 13339 7098 13363 7100
rect 13419 7098 13443 7100
rect 13499 7098 13505 7100
rect 13259 7046 13261 7098
rect 13441 7046 13443 7098
rect 13197 7044 13203 7046
rect 13259 7044 13283 7046
rect 13339 7044 13363 7046
rect 13419 7044 13443 7046
rect 13499 7044 13505 7046
rect 13197 7035 13505 7044
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12360 6322 12388 6938
rect 13832 6934 13860 9046
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 12532 6384 12584 6390
rect 12452 6332 12532 6338
rect 12452 6326 12584 6332
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12452 6310 12572 6326
rect 12452 5642 12480 6310
rect 13197 6012 13505 6021
rect 13197 6010 13203 6012
rect 13259 6010 13283 6012
rect 13339 6010 13363 6012
rect 13419 6010 13443 6012
rect 13499 6010 13505 6012
rect 13259 5958 13261 6010
rect 13441 5958 13443 6010
rect 13197 5956 13203 5958
rect 13259 5956 13283 5958
rect 13339 5956 13363 5958
rect 13419 5956 13443 5958
rect 13499 5956 13505 5958
rect 13197 5947 13505 5956
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12452 5302 12480 5578
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 10747 3292 11055 3301
rect 10747 3290 10753 3292
rect 10809 3290 10833 3292
rect 10889 3290 10913 3292
rect 10969 3290 10993 3292
rect 11049 3290 11055 3292
rect 10809 3238 10811 3290
rect 10991 3238 10993 3290
rect 10747 3236 10753 3238
rect 10809 3236 10833 3238
rect 10889 3236 10913 3238
rect 10969 3236 10993 3238
rect 11049 3236 11055 3238
rect 10747 3227 11055 3236
rect 11348 3126 11376 3402
rect 12452 3126 12480 5238
rect 13832 5234 13860 6870
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13924 5914 13952 6258
rect 14200 6254 14228 10542
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 5370 13952 5646
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 14200 5166 14228 6190
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13197 4924 13505 4933
rect 13197 4922 13203 4924
rect 13259 4922 13283 4924
rect 13339 4922 13363 4924
rect 13419 4922 13443 4924
rect 13499 4922 13505 4924
rect 13259 4870 13261 4922
rect 13441 4870 13443 4922
rect 13197 4868 13203 4870
rect 13259 4868 13283 4870
rect 13339 4868 13363 4870
rect 13419 4868 13443 4870
rect 13499 4868 13505 4870
rect 13197 4859 13505 4868
rect 13197 3836 13505 3845
rect 13197 3834 13203 3836
rect 13259 3834 13283 3836
rect 13339 3834 13363 3836
rect 13419 3834 13443 3836
rect 13499 3834 13505 3836
rect 13259 3782 13261 3834
rect 13441 3782 13443 3834
rect 13197 3780 13203 3782
rect 13259 3780 13283 3782
rect 13339 3780 13363 3782
rect 13419 3780 13443 3782
rect 13499 3780 13505 3782
rect 13197 3771 13505 3780
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2446 11192 2790
rect 12544 2446 12572 3334
rect 13197 2748 13505 2757
rect 13197 2746 13203 2748
rect 13259 2746 13283 2748
rect 13339 2746 13363 2748
rect 13419 2746 13443 2748
rect 13499 2746 13505 2748
rect 13259 2694 13261 2746
rect 13441 2694 13443 2746
rect 13197 2692 13203 2694
rect 13259 2692 13283 2694
rect 13339 2692 13363 2694
rect 13419 2692 13443 2694
rect 13499 2692 13505 2694
rect 13197 2683 13505 2692
rect 14292 2446 14320 10406
rect 14568 9994 14596 12174
rect 14660 10742 14688 12922
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15028 11354 15056 11698
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 15212 10130 15240 11018
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 9994 15240 10066
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15120 8634 15148 8910
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7954 14596 8230
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14568 7410 14596 7890
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15304 6254 15332 6666
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 15028 5914 15056 6122
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 15304 5778 15332 6190
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15304 5534 15332 5714
rect 15212 5506 15332 5534
rect 15212 4690 15240 5506
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15396 4622 15424 6394
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15488 3602 15516 15166
rect 15646 14172 15954 14181
rect 15646 14170 15652 14172
rect 15708 14170 15732 14172
rect 15788 14170 15812 14172
rect 15868 14170 15892 14172
rect 15948 14170 15954 14172
rect 15708 14118 15710 14170
rect 15890 14118 15892 14170
rect 15646 14116 15652 14118
rect 15708 14116 15732 14118
rect 15788 14116 15812 14118
rect 15868 14116 15892 14118
rect 15948 14116 15954 14118
rect 15646 14107 15954 14116
rect 16132 13258 16160 15370
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16500 13326 16528 14894
rect 16592 14618 16620 21490
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 20942 16712 21422
rect 17604 21146 17632 21490
rect 18096 21244 18404 21253
rect 18096 21242 18102 21244
rect 18158 21242 18182 21244
rect 18238 21242 18262 21244
rect 18318 21242 18342 21244
rect 18398 21242 18404 21244
rect 18158 21190 18160 21242
rect 18340 21190 18342 21242
rect 18096 21188 18102 21190
rect 18158 21188 18182 21190
rect 18238 21188 18262 21190
rect 18318 21188 18342 21190
rect 18398 21188 18404 21190
rect 18096 21179 18404 21188
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 18420 20936 18472 20942
rect 18472 20884 18552 20890
rect 18420 20878 18552 20884
rect 17592 20868 17644 20874
rect 18432 20862 18552 20878
rect 17592 20810 17644 20816
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17236 20466 17264 20742
rect 17604 20534 17632 20810
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16776 18086 16804 20334
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17052 18902 17080 19722
rect 17144 19310 17172 19790
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17052 18290 17080 18702
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17236 18222 17264 19110
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17604 18170 17632 20470
rect 17880 19922 17908 20742
rect 18096 20156 18404 20165
rect 18096 20154 18102 20156
rect 18158 20154 18182 20156
rect 18238 20154 18262 20156
rect 18318 20154 18342 20156
rect 18398 20154 18404 20156
rect 18158 20102 18160 20154
rect 18340 20102 18342 20154
rect 18096 20100 18102 20102
rect 18158 20100 18182 20102
rect 18238 20100 18262 20102
rect 18318 20100 18342 20102
rect 18398 20100 18404 20102
rect 18096 20091 18404 20100
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17880 18970 17908 19314
rect 18524 19310 18552 20862
rect 18892 20058 18920 21490
rect 19076 20602 19104 21490
rect 19904 21146 19932 23205
rect 20545 21788 20853 21797
rect 20545 21786 20551 21788
rect 20607 21786 20631 21788
rect 20687 21786 20711 21788
rect 20767 21786 20791 21788
rect 20847 21786 20853 21788
rect 20607 21734 20609 21786
rect 20789 21734 20791 21786
rect 20545 21732 20551 21734
rect 20607 21732 20631 21734
rect 20687 21732 20711 21734
rect 20767 21732 20791 21734
rect 20847 21732 20853 21734
rect 20545 21723 20853 21732
rect 21192 21418 21220 23205
rect 21180 21412 21232 21418
rect 21180 21354 21232 21360
rect 19892 21140 19944 21146
rect 19892 21082 19944 21088
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19260 20602 19288 20946
rect 19892 20936 19944 20942
rect 19430 20904 19486 20913
rect 19892 20878 19944 20884
rect 19430 20839 19486 20848
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19444 20466 19472 20839
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17868 18216 17920 18222
rect 17604 18142 17816 18170
rect 17972 18204 18000 19246
rect 18096 19068 18404 19077
rect 18096 19066 18102 19068
rect 18158 19066 18182 19068
rect 18238 19066 18262 19068
rect 18318 19066 18342 19068
rect 18398 19066 18404 19068
rect 18158 19014 18160 19066
rect 18340 19014 18342 19066
rect 18096 19012 18102 19014
rect 18158 19012 18182 19014
rect 18238 19012 18262 19014
rect 18318 19012 18342 19014
rect 18398 19012 18404 19014
rect 18096 19003 18404 19012
rect 18524 18766 18552 19246
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18156 18358 18184 18566
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17920 18176 18000 18204
rect 17868 18158 17920 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 15646 13084 15954 13093
rect 15646 13082 15652 13084
rect 15708 13082 15732 13084
rect 15788 13082 15812 13084
rect 15868 13082 15892 13084
rect 15948 13082 15954 13084
rect 15708 13030 15710 13082
rect 15890 13030 15892 13082
rect 15646 13028 15652 13030
rect 15708 13028 15732 13030
rect 15788 13028 15812 13030
rect 15868 13028 15892 13030
rect 15948 13028 15954 13030
rect 15646 13019 15954 13028
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 11082 15608 12786
rect 16132 12782 16160 13194
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12170 16160 12718
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 15646 11996 15954 12005
rect 15646 11994 15652 11996
rect 15708 11994 15732 11996
rect 15788 11994 15812 11996
rect 15868 11994 15892 11996
rect 15948 11994 15954 11996
rect 15708 11942 15710 11994
rect 15890 11942 15892 11994
rect 15646 11940 15652 11942
rect 15708 11940 15732 11942
rect 15788 11940 15812 11942
rect 15868 11940 15892 11942
rect 15948 11940 15954 11942
rect 15646 11931 15954 11940
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15856 11354 15884 11562
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15646 10908 15954 10917
rect 15646 10906 15652 10908
rect 15708 10906 15732 10908
rect 15788 10906 15812 10908
rect 15868 10906 15892 10908
rect 15948 10906 15954 10908
rect 15708 10854 15710 10906
rect 15890 10854 15892 10906
rect 15646 10852 15652 10854
rect 15708 10852 15732 10854
rect 15788 10852 15812 10854
rect 15868 10852 15892 10854
rect 15948 10852 15954 10854
rect 15646 10843 15954 10852
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15580 2774 15608 10406
rect 16040 10266 16068 11086
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15646 9820 15954 9829
rect 15646 9818 15652 9820
rect 15708 9818 15732 9820
rect 15788 9818 15812 9820
rect 15868 9818 15892 9820
rect 15948 9818 15954 9820
rect 15708 9766 15710 9818
rect 15890 9766 15892 9818
rect 15646 9764 15652 9766
rect 15708 9764 15732 9766
rect 15788 9764 15812 9766
rect 15868 9764 15892 9766
rect 15948 9764 15954 9766
rect 15646 9755 15954 9764
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15646 8732 15954 8741
rect 15646 8730 15652 8732
rect 15708 8730 15732 8732
rect 15788 8730 15812 8732
rect 15868 8730 15892 8732
rect 15948 8730 15954 8732
rect 15708 8678 15710 8730
rect 15890 8678 15892 8730
rect 15646 8676 15652 8678
rect 15708 8676 15732 8678
rect 15788 8676 15812 8678
rect 15868 8676 15892 8678
rect 15948 8676 15954 8678
rect 15646 8667 15954 8676
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15672 7886 15700 8502
rect 16040 8090 16068 8978
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8566 16160 8774
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16040 7886 16068 8026
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15646 7644 15954 7653
rect 15646 7642 15652 7644
rect 15708 7642 15732 7644
rect 15788 7642 15812 7644
rect 15868 7642 15892 7644
rect 15948 7642 15954 7644
rect 15708 7590 15710 7642
rect 15890 7590 15892 7642
rect 15646 7588 15652 7590
rect 15708 7588 15732 7590
rect 15788 7588 15812 7590
rect 15868 7588 15892 7590
rect 15948 7588 15954 7590
rect 15646 7579 15954 7588
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 6798 15700 7142
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15646 6556 15954 6565
rect 15646 6554 15652 6556
rect 15708 6554 15732 6556
rect 15788 6554 15812 6556
rect 15868 6554 15892 6556
rect 15948 6554 15954 6556
rect 15708 6502 15710 6554
rect 15890 6502 15892 6554
rect 15646 6500 15652 6502
rect 15708 6500 15732 6502
rect 15788 6500 15812 6502
rect 15868 6500 15892 6502
rect 15948 6500 15954 6502
rect 15646 6491 15954 6500
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 15646 5468 15954 5477
rect 15646 5466 15652 5468
rect 15708 5466 15732 5468
rect 15788 5466 15812 5468
rect 15868 5466 15892 5468
rect 15948 5466 15954 5468
rect 15708 5414 15710 5466
rect 15890 5414 15892 5466
rect 15646 5412 15652 5414
rect 15708 5412 15732 5414
rect 15788 5412 15812 5414
rect 15868 5412 15892 5414
rect 15948 5412 15954 5414
rect 15646 5403 15954 5412
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 4758 15976 4966
rect 16040 4826 16068 5782
rect 16132 5166 16160 6122
rect 16224 6118 16252 11222
rect 16592 6390 16620 11698
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15936 4752 15988 4758
rect 16132 4706 16160 5102
rect 15936 4694 15988 4700
rect 16040 4678 16160 4706
rect 15646 4380 15954 4389
rect 15646 4378 15652 4380
rect 15708 4378 15732 4380
rect 15788 4378 15812 4380
rect 15868 4378 15892 4380
rect 15948 4378 15954 4380
rect 15708 4326 15710 4378
rect 15890 4326 15892 4378
rect 15646 4324 15652 4326
rect 15708 4324 15732 4326
rect 15788 4324 15812 4326
rect 15868 4324 15892 4326
rect 15948 4324 15954 4326
rect 15646 4315 15954 4324
rect 16040 3602 16068 4678
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15646 3292 15954 3301
rect 15646 3290 15652 3292
rect 15708 3290 15732 3292
rect 15788 3290 15812 3292
rect 15868 3290 15892 3292
rect 15948 3290 15954 3292
rect 15708 3238 15710 3290
rect 15890 3238 15892 3290
rect 15646 3236 15652 3238
rect 15708 3236 15732 3238
rect 15788 3236 15812 3238
rect 15868 3236 15892 3238
rect 15948 3236 15954 3238
rect 15646 3227 15954 3236
rect 16040 2990 16068 3538
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15396 2746 15608 2774
rect 15396 2446 15424 2746
rect 16684 2446 16712 13126
rect 16776 3058 16804 18022
rect 17788 17746 17816 18142
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17604 17338 17632 17682
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 16658 17540 17070
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17696 16114 17724 17614
rect 17788 17610 17816 17682
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17788 16522 17816 17546
rect 17880 17542 17908 18158
rect 18096 17980 18404 17989
rect 18096 17978 18102 17980
rect 18158 17978 18182 17980
rect 18238 17978 18262 17980
rect 18318 17978 18342 17980
rect 18398 17978 18404 17980
rect 18158 17926 18160 17978
rect 18340 17926 18342 17978
rect 18096 17924 18102 17926
rect 18158 17924 18182 17926
rect 18238 17924 18262 17926
rect 18318 17924 18342 17926
rect 18398 17924 18404 17926
rect 18096 17915 18404 17924
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17202 17908 17478
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 18524 17134 18552 18702
rect 18708 17678 18736 19654
rect 18892 18426 18920 19790
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18984 19446 19012 19722
rect 19444 19514 19472 19858
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18788 18352 18840 18358
rect 18788 18294 18840 18300
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18604 17536 18656 17542
rect 18800 17524 18828 18294
rect 19536 17882 19564 20402
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 18656 17496 18828 17524
rect 18604 17478 18656 17484
rect 18616 17270 18644 17478
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18096 16892 18404 16901
rect 18096 16890 18102 16892
rect 18158 16890 18182 16892
rect 18238 16890 18262 16892
rect 18318 16890 18342 16892
rect 18398 16890 18404 16892
rect 18158 16838 18160 16890
rect 18340 16838 18342 16890
rect 18096 16836 18102 16838
rect 18158 16836 18182 16838
rect 18238 16836 18262 16838
rect 18318 16836 18342 16838
rect 18398 16836 18404 16838
rect 18096 16827 18404 16836
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17788 16182 17816 16458
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 14414 16896 15302
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16960 12986 16988 16050
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18096 15804 18404 15813
rect 18096 15802 18102 15804
rect 18158 15802 18182 15804
rect 18238 15802 18262 15804
rect 18318 15802 18342 15804
rect 18398 15802 18404 15804
rect 18158 15750 18160 15802
rect 18340 15750 18342 15802
rect 18096 15748 18102 15750
rect 18158 15748 18182 15750
rect 18238 15748 18262 15750
rect 18318 15748 18342 15750
rect 18398 15748 18404 15750
rect 18096 15739 18404 15748
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17052 14618 17080 15574
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17420 12442 17448 14486
rect 17604 14482 17632 15506
rect 18432 14958 18460 15982
rect 18524 15502 18552 16390
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 15706 18736 15982
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15094 18736 15302
rect 19352 15094 19380 15370
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18096 14716 18404 14725
rect 18096 14714 18102 14716
rect 18158 14714 18182 14716
rect 18238 14714 18262 14716
rect 18318 14714 18342 14716
rect 18398 14714 18404 14716
rect 18158 14662 18160 14714
rect 18340 14662 18342 14714
rect 18096 14660 18102 14662
rect 18158 14660 18182 14662
rect 18238 14660 18262 14662
rect 18318 14660 18342 14662
rect 18398 14660 18404 14662
rect 18096 14651 18404 14660
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 14006 18460 14214
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18800 13870 18828 14894
rect 19352 14006 19380 15030
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18096 13628 18404 13637
rect 18096 13626 18102 13628
rect 18158 13626 18182 13628
rect 18238 13626 18262 13628
rect 18318 13626 18342 13628
rect 18398 13626 18404 13628
rect 18158 13574 18160 13626
rect 18340 13574 18342 13626
rect 18096 13572 18102 13574
rect 18158 13572 18182 13574
rect 18238 13572 18262 13574
rect 18318 13572 18342 13574
rect 18398 13572 18404 13574
rect 18096 13563 18404 13572
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16960 11762 16988 12038
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16856 11688 16908 11694
rect 16908 11636 16988 11642
rect 16856 11630 16988 11636
rect 16868 11614 16988 11630
rect 16960 11218 16988 11614
rect 17788 11354 17816 12718
rect 18096 12540 18404 12549
rect 18096 12538 18102 12540
rect 18158 12538 18182 12540
rect 18238 12538 18262 12540
rect 18318 12538 18342 12540
rect 18398 12538 18404 12540
rect 18158 12486 18160 12538
rect 18340 12486 18342 12538
rect 18096 12484 18102 12486
rect 18158 12484 18182 12486
rect 18238 12484 18262 12486
rect 18318 12484 18342 12486
rect 18398 12484 18404 12486
rect 18096 12475 18404 12484
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18064 11694 18092 12242
rect 18156 11898 18184 12310
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18052 11688 18104 11694
rect 17972 11636 18052 11642
rect 17972 11630 18104 11636
rect 17972 11614 18092 11630
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17972 11218 18000 11614
rect 18096 11452 18404 11461
rect 18096 11450 18102 11452
rect 18158 11450 18182 11452
rect 18238 11450 18262 11452
rect 18318 11450 18342 11452
rect 18398 11450 18404 11452
rect 18158 11398 18160 11450
rect 18340 11398 18342 11450
rect 18096 11396 18102 11398
rect 18158 11396 18182 11398
rect 18238 11396 18262 11398
rect 18318 11396 18342 11398
rect 18398 11396 18404 11398
rect 18096 11387 18404 11396
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 9654 17264 10950
rect 17880 10810 17908 11086
rect 18432 11054 18460 12718
rect 18616 12238 18644 13126
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18708 12442 18736 12718
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18432 11026 18552 11054
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17788 9722 17816 10610
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18096 10364 18404 10373
rect 18096 10362 18102 10364
rect 18158 10362 18182 10364
rect 18238 10362 18262 10364
rect 18318 10362 18342 10364
rect 18398 10362 18404 10364
rect 18158 10310 18160 10362
rect 18340 10310 18342 10362
rect 18096 10308 18102 10310
rect 18158 10308 18182 10310
rect 18238 10308 18262 10310
rect 18318 10308 18342 10310
rect 18398 10308 18404 10310
rect 18096 10299 18404 10308
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17880 9110 17908 9454
rect 17972 9178 18000 9522
rect 18432 9518 18460 10542
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18096 9276 18404 9285
rect 18096 9274 18102 9276
rect 18158 9274 18182 9276
rect 18238 9274 18262 9276
rect 18318 9274 18342 9276
rect 18398 9274 18404 9276
rect 18158 9222 18160 9274
rect 18340 9222 18342 9274
rect 18096 9220 18102 9222
rect 18158 9220 18182 9222
rect 18238 9220 18262 9222
rect 18318 9220 18342 9222
rect 18398 9220 18404 9222
rect 18096 9211 18404 9220
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8566 17172 8910
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17604 8566 17632 8842
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 7410 17816 8230
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17880 7342 17908 9046
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18096 8188 18404 8197
rect 18096 8186 18102 8188
rect 18158 8186 18182 8188
rect 18238 8186 18262 8188
rect 18318 8186 18342 8188
rect 18398 8186 18404 8188
rect 18158 8134 18160 8186
rect 18340 8134 18342 8186
rect 18096 8132 18102 8134
rect 18158 8132 18182 8134
rect 18238 8132 18262 8134
rect 18318 8132 18342 8134
rect 18398 8132 18404 8134
rect 18096 8123 18404 8132
rect 18432 8022 18460 8910
rect 18524 8090 18552 11026
rect 18708 10742 18736 11494
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18800 10606 18828 13806
rect 19352 12918 19380 13942
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19352 10742 19380 12854
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 19352 9654 19380 10678
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19352 8906 19380 9590
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8498 19288 8774
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 19076 7886 19104 8230
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19352 7478 19380 8842
rect 19628 8090 19656 8842
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19628 7546 19656 7822
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 6322 16896 6598
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17052 5534 17080 6326
rect 17144 5710 17172 7278
rect 18096 7100 18404 7109
rect 18096 7098 18102 7100
rect 18158 7098 18182 7100
rect 18238 7098 18262 7100
rect 18318 7098 18342 7100
rect 18398 7098 18404 7100
rect 18158 7046 18160 7098
rect 18340 7046 18342 7098
rect 18096 7044 18102 7046
rect 18158 7044 18182 7046
rect 18238 7044 18262 7046
rect 18318 7044 18342 7046
rect 18398 7044 18404 7046
rect 18096 7035 18404 7044
rect 18708 6458 18736 7278
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18096 6012 18404 6021
rect 18096 6010 18102 6012
rect 18158 6010 18182 6012
rect 18238 6010 18262 6012
rect 18318 6010 18342 6012
rect 18398 6010 18404 6012
rect 18158 5958 18160 6010
rect 18340 5958 18342 6010
rect 18096 5956 18102 5958
rect 18158 5956 18182 5958
rect 18238 5956 18262 5958
rect 18318 5956 18342 5958
rect 18398 5956 18404 5958
rect 18096 5947 18404 5956
rect 18616 5778 18644 6054
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 16960 5506 17080 5534
rect 16960 5302 16988 5506
rect 16948 5296 17000 5302
rect 16868 5244 16948 5250
rect 16868 5238 17000 5244
rect 16868 5222 16988 5238
rect 17144 5234 17172 5646
rect 19352 5642 19380 7414
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 17512 5302 17540 5510
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 17132 5228 17184 5234
rect 16868 3466 16896 5222
rect 17132 5170 17184 5176
rect 17144 4146 17172 5170
rect 18096 4924 18404 4933
rect 18096 4922 18102 4924
rect 18158 4922 18182 4924
rect 18238 4922 18262 4924
rect 18318 4922 18342 4924
rect 18398 4922 18404 4924
rect 18158 4870 18160 4922
rect 18340 4870 18342 4922
rect 18096 4868 18102 4870
rect 18158 4868 18182 4870
rect 18238 4868 18262 4870
rect 18318 4868 18342 4870
rect 18398 4868 18404 4870
rect 18096 4859 18404 4868
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17696 4010 17724 4422
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 18096 3836 18404 3845
rect 18096 3834 18102 3836
rect 18158 3834 18182 3836
rect 18238 3834 18262 3836
rect 18318 3834 18342 3836
rect 18398 3834 18404 3836
rect 18158 3782 18160 3834
rect 18340 3782 18342 3834
rect 18096 3780 18102 3782
rect 18158 3780 18182 3782
rect 18238 3780 18262 3782
rect 18318 3780 18342 3782
rect 18398 3780 18404 3782
rect 18096 3771 18404 3780
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 3194 16896 3402
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 17420 2446 17448 3334
rect 18892 3058 18920 5510
rect 19352 5302 19380 5578
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19352 4214 19380 5238
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 18096 2748 18404 2757
rect 18096 2746 18102 2748
rect 18158 2746 18182 2748
rect 18238 2746 18262 2748
rect 18318 2746 18342 2748
rect 18398 2746 18404 2748
rect 18158 2694 18160 2746
rect 18340 2694 18342 2746
rect 18096 2692 18102 2694
rect 18158 2692 18182 2694
rect 18238 2692 18262 2694
rect 18318 2692 18342 2694
rect 18398 2692 18404 2694
rect 18096 2683 18404 2692
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 5848 2204 6156 2213
rect 5848 2202 5854 2204
rect 5910 2202 5934 2204
rect 5990 2202 6014 2204
rect 6070 2202 6094 2204
rect 6150 2202 6156 2204
rect 5910 2150 5912 2202
rect 6092 2150 6094 2202
rect 5848 2148 5854 2150
rect 5910 2148 5934 2150
rect 5990 2148 6014 2150
rect 6070 2148 6094 2150
rect 6150 2148 6156 2150
rect 5848 2139 6156 2148
rect 7024 800 7052 2246
rect 8312 800 8340 2246
rect 9600 800 9628 2246
rect 570 0 626 800
rect 1858 0 1914 800
rect 3146 0 3202 800
rect 4434 0 4490 800
rect 5722 0 5778 800
rect 7010 0 7066 800
rect 8298 0 8354 800
rect 9586 0 9642 800
rect 10612 762 10640 2246
rect 10747 2204 11055 2213
rect 10747 2202 10753 2204
rect 10809 2202 10833 2204
rect 10889 2202 10913 2204
rect 10969 2202 10993 2204
rect 11049 2202 11055 2204
rect 10809 2150 10811 2202
rect 10991 2150 10993 2202
rect 10747 2148 10753 2150
rect 10809 2148 10833 2150
rect 10889 2148 10913 2150
rect 10969 2148 10993 2150
rect 11049 2148 11055 2150
rect 10747 2139 11055 2148
rect 10796 870 10916 898
rect 10796 762 10824 870
rect 10888 800 10916 870
rect 12176 800 12204 2246
rect 13464 800 13492 2246
rect 14752 800 14780 2246
rect 15646 2204 15954 2213
rect 15646 2202 15652 2204
rect 15708 2202 15732 2204
rect 15788 2202 15812 2204
rect 15868 2202 15892 2204
rect 15948 2202 15954 2204
rect 15708 2150 15710 2202
rect 15890 2150 15892 2202
rect 15646 2148 15652 2150
rect 15708 2148 15732 2150
rect 15788 2148 15812 2150
rect 15868 2148 15892 2150
rect 15948 2148 15954 2150
rect 15646 2139 15954 2148
rect 16040 800 16068 2246
rect 17328 800 17356 2246
rect 18616 870 18736 898
rect 18616 800 18644 870
rect 10612 734 10824 762
rect 10874 0 10930 800
rect 12162 0 12218 800
rect 13450 0 13506 800
rect 14738 0 14794 800
rect 16026 0 16082 800
rect 17314 0 17370 800
rect 18602 0 18658 800
rect 18708 762 18736 870
rect 18892 762 18920 2246
rect 19168 1465 19196 2790
rect 19260 2650 19288 2858
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19444 2446 19472 2926
rect 19720 2514 19748 19110
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19812 17610 19840 18838
rect 19904 18426 19932 20878
rect 20545 20700 20853 20709
rect 20545 20698 20551 20700
rect 20607 20698 20631 20700
rect 20687 20698 20711 20700
rect 20767 20698 20791 20700
rect 20847 20698 20853 20700
rect 20607 20646 20609 20698
rect 20789 20646 20791 20698
rect 20545 20644 20551 20646
rect 20607 20644 20631 20646
rect 20687 20644 20711 20646
rect 20767 20644 20791 20646
rect 20847 20644 20853 20646
rect 20545 20635 20853 20644
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20088 19145 20116 20198
rect 20545 19612 20853 19621
rect 20545 19610 20551 19612
rect 20607 19610 20631 19612
rect 20687 19610 20711 19612
rect 20767 19610 20791 19612
rect 20847 19610 20853 19612
rect 20607 19558 20609 19610
rect 20789 19558 20791 19610
rect 20545 19556 20551 19558
rect 20607 19556 20631 19558
rect 20687 19556 20711 19558
rect 20767 19556 20791 19558
rect 20847 19556 20853 19558
rect 20545 19547 20853 19556
rect 20074 19136 20130 19145
rect 20074 19071 20130 19080
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19996 17921 20024 18566
rect 19982 17912 20038 17921
rect 19982 17847 20038 17856
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19812 16114 19840 17546
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19904 5534 19932 16934
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 15609 20024 16390
rect 19982 15600 20038 15609
rect 19982 15535 20038 15544
rect 20088 15502 20116 17546
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20180 15162 20208 16526
rect 20272 16250 20300 18702
rect 20545 18524 20853 18533
rect 20545 18522 20551 18524
rect 20607 18522 20631 18524
rect 20687 18522 20711 18524
rect 20767 18522 20791 18524
rect 20847 18522 20853 18524
rect 20607 18470 20609 18522
rect 20789 18470 20791 18522
rect 20545 18468 20551 18470
rect 20607 18468 20631 18470
rect 20687 18468 20711 18470
rect 20767 18468 20791 18470
rect 20847 18468 20853 18470
rect 20545 18459 20853 18468
rect 20545 17436 20853 17445
rect 20545 17434 20551 17436
rect 20607 17434 20631 17436
rect 20687 17434 20711 17436
rect 20767 17434 20791 17436
rect 20847 17434 20853 17436
rect 20607 17382 20609 17434
rect 20789 17382 20791 17434
rect 20545 17380 20551 17382
rect 20607 17380 20631 17382
rect 20687 17380 20711 17382
rect 20767 17380 20791 17382
rect 20847 17380 20853 17382
rect 20545 17371 20853 17380
rect 20545 16348 20853 16357
rect 20545 16346 20551 16348
rect 20607 16346 20631 16348
rect 20687 16346 20711 16348
rect 20767 16346 20791 16348
rect 20847 16346 20853 16348
rect 20607 16294 20609 16346
rect 20789 16294 20791 16346
rect 20545 16292 20551 16294
rect 20607 16292 20631 16294
rect 20687 16292 20711 16294
rect 20767 16292 20791 16294
rect 20847 16292 20853 16294
rect 20545 16283 20853 16292
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20545 15260 20853 15269
rect 20545 15258 20551 15260
rect 20607 15258 20631 15260
rect 20687 15258 20711 15260
rect 20767 15258 20791 15260
rect 20847 15258 20853 15260
rect 20607 15206 20609 15258
rect 20789 15206 20791 15258
rect 20545 15204 20551 15206
rect 20607 15204 20631 15206
rect 20687 15204 20711 15206
rect 20767 15204 20791 15206
rect 20847 15204 20853 15206
rect 20545 15195 20853 15204
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20545 14172 20853 14181
rect 20545 14170 20551 14172
rect 20607 14170 20631 14172
rect 20687 14170 20711 14172
rect 20767 14170 20791 14172
rect 20847 14170 20853 14172
rect 20607 14118 20609 14170
rect 20789 14118 20791 14170
rect 20545 14116 20551 14118
rect 20607 14116 20631 14118
rect 20687 14116 20711 14118
rect 20767 14116 20791 14118
rect 20847 14116 20853 14118
rect 20545 14107 20853 14116
rect 19982 13832 20038 13841
rect 19982 13767 20038 13776
rect 19996 13530 20024 13767
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20180 13326 20208 13670
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20545 13084 20853 13093
rect 20545 13082 20551 13084
rect 20607 13082 20631 13084
rect 20687 13082 20711 13084
rect 20767 13082 20791 13084
rect 20847 13082 20853 13084
rect 20607 13030 20609 13082
rect 20789 13030 20791 13082
rect 20545 13028 20551 13030
rect 20607 13028 20631 13030
rect 20687 13028 20711 13030
rect 20767 13028 20791 13030
rect 20847 13028 20853 13030
rect 20545 13019 20853 13028
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 19984 12368 20036 12374
rect 19982 12336 19984 12345
rect 20036 12336 20038 12345
rect 19982 12271 20038 12280
rect 20180 12238 20208 12582
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20545 11996 20853 12005
rect 20545 11994 20551 11996
rect 20607 11994 20631 11996
rect 20687 11994 20711 11996
rect 20767 11994 20791 11996
rect 20847 11994 20853 11996
rect 20607 11942 20609 11994
rect 20789 11942 20791 11994
rect 20545 11940 20551 11942
rect 20607 11940 20631 11942
rect 20687 11940 20711 11942
rect 20767 11940 20791 11942
rect 20847 11940 20853 11942
rect 20545 11931 20853 11940
rect 20545 10908 20853 10917
rect 20545 10906 20551 10908
rect 20607 10906 20631 10908
rect 20687 10906 20711 10908
rect 20767 10906 20791 10908
rect 20847 10906 20853 10908
rect 20607 10854 20609 10906
rect 20789 10854 20791 10906
rect 20545 10852 20551 10854
rect 20607 10852 20631 10854
rect 20687 10852 20711 10854
rect 20767 10852 20791 10854
rect 20847 10852 20853 10854
rect 20545 10843 20853 10852
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19982 10296 20038 10305
rect 19982 10231 19984 10240
rect 20036 10231 20038 10240
rect 19984 10202 20036 10208
rect 20180 10062 20208 10406
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20545 9820 20853 9829
rect 20545 9818 20551 9820
rect 20607 9818 20631 9820
rect 20687 9818 20711 9820
rect 20767 9818 20791 9820
rect 20847 9818 20853 9820
rect 20607 9766 20609 9818
rect 20789 9766 20791 9818
rect 20545 9764 20551 9766
rect 20607 9764 20631 9766
rect 20687 9764 20711 9766
rect 20767 9764 20791 9766
rect 20847 9764 20853 9766
rect 20545 9755 20853 9764
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19996 8537 20024 8570
rect 19982 8528 20038 8537
rect 20180 8498 20208 9318
rect 20545 8732 20853 8741
rect 20545 8730 20551 8732
rect 20607 8730 20631 8732
rect 20687 8730 20711 8732
rect 20767 8730 20791 8732
rect 20847 8730 20853 8732
rect 20607 8678 20609 8730
rect 20789 8678 20791 8730
rect 20545 8676 20551 8678
rect 20607 8676 20631 8678
rect 20687 8676 20711 8678
rect 20767 8676 20791 8678
rect 20847 8676 20853 8678
rect 20545 8667 20853 8676
rect 19982 8463 20038 8472
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20545 7644 20853 7653
rect 20545 7642 20551 7644
rect 20607 7642 20631 7644
rect 20687 7642 20711 7644
rect 20767 7642 20791 7644
rect 20847 7642 20853 7644
rect 20607 7590 20609 7642
rect 20789 7590 20791 7642
rect 20545 7588 20551 7590
rect 20607 7588 20631 7590
rect 20687 7588 20711 7590
rect 20767 7588 20791 7590
rect 20847 7588 20853 7590
rect 20545 7579 20853 7588
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20180 6798 20208 7142
rect 20168 6792 20220 6798
rect 19982 6760 20038 6769
rect 20168 6734 20220 6740
rect 19982 6695 20038 6704
rect 19996 6662 20024 6695
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 20545 6556 20853 6565
rect 20545 6554 20551 6556
rect 20607 6554 20631 6556
rect 20687 6554 20711 6556
rect 20767 6554 20791 6556
rect 20847 6554 20853 6556
rect 20607 6502 20609 6554
rect 20789 6502 20791 6554
rect 20545 6500 20551 6502
rect 20607 6500 20631 6502
rect 20687 6500 20711 6502
rect 20767 6500 20791 6502
rect 20847 6500 20853 6502
rect 20545 6491 20853 6500
rect 19812 5506 19932 5534
rect 19812 3058 19840 5506
rect 20545 5468 20853 5477
rect 20545 5466 20551 5468
rect 20607 5466 20631 5468
rect 20687 5466 20711 5468
rect 20767 5466 20791 5468
rect 20847 5466 20853 5468
rect 20607 5414 20609 5466
rect 20789 5414 20791 5466
rect 20545 5412 20551 5414
rect 20607 5412 20631 5414
rect 20687 5412 20711 5414
rect 20767 5412 20791 5414
rect 20847 5412 20853 5414
rect 20545 5403 20853 5412
rect 20076 5024 20128 5030
rect 20074 4992 20076 5001
rect 20128 4992 20130 5001
rect 20074 4927 20130 4936
rect 20545 4380 20853 4389
rect 20545 4378 20551 4380
rect 20607 4378 20631 4380
rect 20687 4378 20711 4380
rect 20767 4378 20791 4380
rect 20847 4378 20853 4380
rect 20607 4326 20609 4378
rect 20789 4326 20791 4378
rect 20545 4324 20551 4326
rect 20607 4324 20631 4326
rect 20687 4324 20711 4326
rect 20767 4324 20791 4326
rect 20847 4324 20853 4326
rect 20545 4315 20853 4324
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19904 3534 19932 3878
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 20074 3496 20130 3505
rect 20074 3431 20130 3440
rect 20088 3398 20116 3431
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20545 3292 20853 3301
rect 20545 3290 20551 3292
rect 20607 3290 20631 3292
rect 20687 3290 20711 3292
rect 20767 3290 20791 3292
rect 20847 3290 20853 3292
rect 20607 3238 20609 3290
rect 20789 3238 20791 3290
rect 20545 3236 20551 3238
rect 20607 3236 20631 3238
rect 20687 3236 20711 3238
rect 20767 3236 20791 3238
rect 20847 3236 20853 3238
rect 20545 3227 20853 3236
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 21180 2916 21232 2922
rect 21180 2858 21232 2864
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19154 1456 19210 1465
rect 19154 1391 19210 1400
rect 19904 800 19932 2790
rect 20545 2204 20853 2213
rect 20545 2202 20551 2204
rect 20607 2202 20631 2204
rect 20687 2202 20711 2204
rect 20767 2202 20791 2204
rect 20847 2202 20853 2204
rect 20607 2150 20609 2202
rect 20789 2150 20791 2202
rect 20545 2148 20551 2150
rect 20607 2148 20631 2150
rect 20687 2148 20711 2150
rect 20767 2148 20791 2150
rect 20847 2148 20853 2150
rect 20545 2139 20853 2148
rect 21192 800 21220 2858
rect 18708 734 18920 762
rect 19890 0 19946 800
rect 21178 0 21234 800
<< via2 >>
rect 1674 21800 1730 21856
rect 1120 18460 1470 18540
rect 5854 21786 5910 21788
rect 5934 21786 5990 21788
rect 6014 21786 6070 21788
rect 6094 21786 6150 21788
rect 5854 21734 5900 21786
rect 5900 21734 5910 21786
rect 5934 21734 5964 21786
rect 5964 21734 5976 21786
rect 5976 21734 5990 21786
rect 6014 21734 6028 21786
rect 6028 21734 6040 21786
rect 6040 21734 6070 21786
rect 6094 21734 6104 21786
rect 6104 21734 6150 21786
rect 5854 21732 5910 21734
rect 5934 21732 5990 21734
rect 6014 21732 6070 21734
rect 6094 21732 6150 21734
rect 10753 21786 10809 21788
rect 10833 21786 10889 21788
rect 10913 21786 10969 21788
rect 10993 21786 11049 21788
rect 10753 21734 10799 21786
rect 10799 21734 10809 21786
rect 10833 21734 10863 21786
rect 10863 21734 10875 21786
rect 10875 21734 10889 21786
rect 10913 21734 10927 21786
rect 10927 21734 10939 21786
rect 10939 21734 10969 21786
rect 10993 21734 11003 21786
rect 11003 21734 11049 21786
rect 10753 21732 10809 21734
rect 10833 21732 10889 21734
rect 10913 21732 10969 21734
rect 10993 21732 11049 21734
rect 15652 21786 15708 21788
rect 15732 21786 15788 21788
rect 15812 21786 15868 21788
rect 15892 21786 15948 21788
rect 15652 21734 15698 21786
rect 15698 21734 15708 21786
rect 15732 21734 15762 21786
rect 15762 21734 15774 21786
rect 15774 21734 15788 21786
rect 15812 21734 15826 21786
rect 15826 21734 15838 21786
rect 15838 21734 15868 21786
rect 15892 21734 15902 21786
rect 15902 21734 15948 21786
rect 15652 21732 15708 21734
rect 15732 21732 15788 21734
rect 15812 21732 15868 21734
rect 15892 21732 15948 21734
rect 16486 22616 16542 22672
rect 1582 13912 1638 13968
rect 1582 9968 1638 10024
rect 3405 21242 3461 21244
rect 3485 21242 3541 21244
rect 3565 21242 3621 21244
rect 3645 21242 3701 21244
rect 3405 21190 3451 21242
rect 3451 21190 3461 21242
rect 3485 21190 3515 21242
rect 3515 21190 3527 21242
rect 3527 21190 3541 21242
rect 3565 21190 3579 21242
rect 3579 21190 3591 21242
rect 3591 21190 3621 21242
rect 3645 21190 3655 21242
rect 3655 21190 3701 21242
rect 3405 21188 3461 21190
rect 3485 21188 3541 21190
rect 3565 21188 3621 21190
rect 3645 21188 3701 21190
rect 3405 20154 3461 20156
rect 3485 20154 3541 20156
rect 3565 20154 3621 20156
rect 3645 20154 3701 20156
rect 3405 20102 3451 20154
rect 3451 20102 3461 20154
rect 3485 20102 3515 20154
rect 3515 20102 3527 20154
rect 3527 20102 3541 20154
rect 3565 20102 3579 20154
rect 3579 20102 3591 20154
rect 3591 20102 3621 20154
rect 3645 20102 3655 20154
rect 3655 20102 3701 20154
rect 3405 20100 3461 20102
rect 3485 20100 3541 20102
rect 3565 20100 3621 20102
rect 3645 20100 3701 20102
rect 3405 19066 3461 19068
rect 3485 19066 3541 19068
rect 3565 19066 3621 19068
rect 3645 19066 3701 19068
rect 3405 19014 3451 19066
rect 3451 19014 3461 19066
rect 3485 19014 3515 19066
rect 3515 19014 3527 19066
rect 3527 19014 3541 19066
rect 3565 19014 3579 19066
rect 3579 19014 3591 19066
rect 3591 19014 3621 19066
rect 3645 19014 3655 19066
rect 3655 19014 3701 19066
rect 3405 19012 3461 19014
rect 3485 19012 3541 19014
rect 3565 19012 3621 19014
rect 3645 19012 3701 19014
rect 3405 17978 3461 17980
rect 3485 17978 3541 17980
rect 3565 17978 3621 17980
rect 3645 17978 3701 17980
rect 3405 17926 3451 17978
rect 3451 17926 3461 17978
rect 3485 17926 3515 17978
rect 3515 17926 3527 17978
rect 3527 17926 3541 17978
rect 3565 17926 3579 17978
rect 3579 17926 3591 17978
rect 3591 17926 3621 17978
rect 3645 17926 3655 17978
rect 3655 17926 3701 17978
rect 3405 17924 3461 17926
rect 3485 17924 3541 17926
rect 3565 17924 3621 17926
rect 3645 17924 3701 17926
rect 3405 16890 3461 16892
rect 3485 16890 3541 16892
rect 3565 16890 3621 16892
rect 3645 16890 3701 16892
rect 3405 16838 3451 16890
rect 3451 16838 3461 16890
rect 3485 16838 3515 16890
rect 3515 16838 3527 16890
rect 3527 16838 3541 16890
rect 3565 16838 3579 16890
rect 3579 16838 3591 16890
rect 3591 16838 3621 16890
rect 3645 16838 3655 16890
rect 3655 16838 3701 16890
rect 3405 16836 3461 16838
rect 3485 16836 3541 16838
rect 3565 16836 3621 16838
rect 3645 16836 3701 16838
rect 3405 15802 3461 15804
rect 3485 15802 3541 15804
rect 3565 15802 3621 15804
rect 3645 15802 3701 15804
rect 3405 15750 3451 15802
rect 3451 15750 3461 15802
rect 3485 15750 3515 15802
rect 3515 15750 3527 15802
rect 3527 15750 3541 15802
rect 3565 15750 3579 15802
rect 3579 15750 3591 15802
rect 3591 15750 3621 15802
rect 3645 15750 3655 15802
rect 3655 15750 3701 15802
rect 3405 15748 3461 15750
rect 3485 15748 3541 15750
rect 3565 15748 3621 15750
rect 3645 15748 3701 15750
rect 3405 14714 3461 14716
rect 3485 14714 3541 14716
rect 3565 14714 3621 14716
rect 3645 14714 3701 14716
rect 3405 14662 3451 14714
rect 3451 14662 3461 14714
rect 3485 14662 3515 14714
rect 3515 14662 3527 14714
rect 3527 14662 3541 14714
rect 3565 14662 3579 14714
rect 3579 14662 3591 14714
rect 3591 14662 3621 14714
rect 3645 14662 3655 14714
rect 3655 14662 3701 14714
rect 3405 14660 3461 14662
rect 3485 14660 3541 14662
rect 3565 14660 3621 14662
rect 3645 14660 3701 14662
rect 3405 13626 3461 13628
rect 3485 13626 3541 13628
rect 3565 13626 3621 13628
rect 3645 13626 3701 13628
rect 3405 13574 3451 13626
rect 3451 13574 3461 13626
rect 3485 13574 3515 13626
rect 3515 13574 3527 13626
rect 3527 13574 3541 13626
rect 3565 13574 3579 13626
rect 3579 13574 3591 13626
rect 3591 13574 3621 13626
rect 3645 13574 3655 13626
rect 3655 13574 3701 13626
rect 3405 13572 3461 13574
rect 3485 13572 3541 13574
rect 3565 13572 3621 13574
rect 3645 13572 3701 13574
rect 3405 12538 3461 12540
rect 3485 12538 3541 12540
rect 3565 12538 3621 12540
rect 3645 12538 3701 12540
rect 3405 12486 3451 12538
rect 3451 12486 3461 12538
rect 3485 12486 3515 12538
rect 3515 12486 3527 12538
rect 3527 12486 3541 12538
rect 3565 12486 3579 12538
rect 3579 12486 3591 12538
rect 3591 12486 3621 12538
rect 3645 12486 3655 12538
rect 3655 12486 3701 12538
rect 3405 12484 3461 12486
rect 3485 12484 3541 12486
rect 3565 12484 3621 12486
rect 3645 12484 3701 12486
rect 3405 11450 3461 11452
rect 3485 11450 3541 11452
rect 3565 11450 3621 11452
rect 3645 11450 3701 11452
rect 3405 11398 3451 11450
rect 3451 11398 3461 11450
rect 3485 11398 3515 11450
rect 3515 11398 3527 11450
rect 3527 11398 3541 11450
rect 3565 11398 3579 11450
rect 3579 11398 3591 11450
rect 3591 11398 3621 11450
rect 3645 11398 3655 11450
rect 3655 11398 3701 11450
rect 3405 11396 3461 11398
rect 3485 11396 3541 11398
rect 3565 11396 3621 11398
rect 3645 11396 3701 11398
rect 3405 10362 3461 10364
rect 3485 10362 3541 10364
rect 3565 10362 3621 10364
rect 3645 10362 3701 10364
rect 3405 10310 3451 10362
rect 3451 10310 3461 10362
rect 3485 10310 3515 10362
rect 3515 10310 3527 10362
rect 3527 10310 3541 10362
rect 3565 10310 3579 10362
rect 3579 10310 3591 10362
rect 3591 10310 3621 10362
rect 3645 10310 3655 10362
rect 3655 10310 3701 10362
rect 3405 10308 3461 10310
rect 3485 10308 3541 10310
rect 3565 10308 3621 10310
rect 3645 10308 3701 10310
rect 5854 20698 5910 20700
rect 5934 20698 5990 20700
rect 6014 20698 6070 20700
rect 6094 20698 6150 20700
rect 5854 20646 5900 20698
rect 5900 20646 5910 20698
rect 5934 20646 5964 20698
rect 5964 20646 5976 20698
rect 5976 20646 5990 20698
rect 6014 20646 6028 20698
rect 6028 20646 6040 20698
rect 6040 20646 6070 20698
rect 6094 20646 6104 20698
rect 6104 20646 6150 20698
rect 5854 20644 5910 20646
rect 5934 20644 5990 20646
rect 6014 20644 6070 20646
rect 6094 20644 6150 20646
rect 5854 19610 5910 19612
rect 5934 19610 5990 19612
rect 6014 19610 6070 19612
rect 6094 19610 6150 19612
rect 5854 19558 5900 19610
rect 5900 19558 5910 19610
rect 5934 19558 5964 19610
rect 5964 19558 5976 19610
rect 5976 19558 5990 19610
rect 6014 19558 6028 19610
rect 6028 19558 6040 19610
rect 6040 19558 6070 19610
rect 6094 19558 6104 19610
rect 6104 19558 6150 19610
rect 5854 19556 5910 19558
rect 5934 19556 5990 19558
rect 6014 19556 6070 19558
rect 6094 19556 6150 19558
rect 3405 9274 3461 9276
rect 3485 9274 3541 9276
rect 3565 9274 3621 9276
rect 3645 9274 3701 9276
rect 3405 9222 3451 9274
rect 3451 9222 3461 9274
rect 3485 9222 3515 9274
rect 3515 9222 3527 9274
rect 3527 9222 3541 9274
rect 3565 9222 3579 9274
rect 3579 9222 3591 9274
rect 3591 9222 3621 9274
rect 3645 9222 3655 9274
rect 3655 9222 3701 9274
rect 3405 9220 3461 9222
rect 3485 9220 3541 9222
rect 3565 9220 3621 9222
rect 3645 9220 3701 9222
rect 3405 8186 3461 8188
rect 3485 8186 3541 8188
rect 3565 8186 3621 8188
rect 3645 8186 3701 8188
rect 3405 8134 3451 8186
rect 3451 8134 3461 8186
rect 3485 8134 3515 8186
rect 3515 8134 3527 8186
rect 3527 8134 3541 8186
rect 3565 8134 3579 8186
rect 3579 8134 3591 8186
rect 3591 8134 3621 8186
rect 3645 8134 3655 8186
rect 3655 8134 3701 8186
rect 3405 8132 3461 8134
rect 3485 8132 3541 8134
rect 3565 8132 3621 8134
rect 3645 8132 3701 8134
rect 3405 7098 3461 7100
rect 3485 7098 3541 7100
rect 3565 7098 3621 7100
rect 3645 7098 3701 7100
rect 3405 7046 3451 7098
rect 3451 7046 3461 7098
rect 3485 7046 3515 7098
rect 3515 7046 3527 7098
rect 3527 7046 3541 7098
rect 3565 7046 3579 7098
rect 3579 7046 3591 7098
rect 3591 7046 3621 7098
rect 3645 7046 3655 7098
rect 3655 7046 3701 7098
rect 3405 7044 3461 7046
rect 3485 7044 3541 7046
rect 3565 7044 3621 7046
rect 3645 7044 3701 7046
rect 3405 6010 3461 6012
rect 3485 6010 3541 6012
rect 3565 6010 3621 6012
rect 3645 6010 3701 6012
rect 3405 5958 3451 6010
rect 3451 5958 3461 6010
rect 3485 5958 3515 6010
rect 3515 5958 3527 6010
rect 3527 5958 3541 6010
rect 3565 5958 3579 6010
rect 3579 5958 3591 6010
rect 3591 5958 3621 6010
rect 3645 5958 3655 6010
rect 3655 5958 3701 6010
rect 3405 5956 3461 5958
rect 3485 5956 3541 5958
rect 3565 5956 3621 5958
rect 3645 5956 3701 5958
rect 3405 4922 3461 4924
rect 3485 4922 3541 4924
rect 3565 4922 3621 4924
rect 3645 4922 3701 4924
rect 3405 4870 3451 4922
rect 3451 4870 3461 4922
rect 3485 4870 3515 4922
rect 3515 4870 3527 4922
rect 3527 4870 3541 4922
rect 3565 4870 3579 4922
rect 3579 4870 3591 4922
rect 3591 4870 3621 4922
rect 3645 4870 3655 4922
rect 3655 4870 3701 4922
rect 3405 4868 3461 4870
rect 3485 4868 3541 4870
rect 3565 4868 3621 4870
rect 3645 4868 3701 4870
rect 1766 2080 1822 2136
rect 3405 3834 3461 3836
rect 3485 3834 3541 3836
rect 3565 3834 3621 3836
rect 3645 3834 3701 3836
rect 3405 3782 3451 3834
rect 3451 3782 3461 3834
rect 3485 3782 3515 3834
rect 3515 3782 3527 3834
rect 3527 3782 3541 3834
rect 3565 3782 3579 3834
rect 3579 3782 3591 3834
rect 3591 3782 3621 3834
rect 3645 3782 3655 3834
rect 3655 3782 3701 3834
rect 3405 3780 3461 3782
rect 3485 3780 3541 3782
rect 3565 3780 3621 3782
rect 3645 3780 3701 3782
rect 3405 2746 3461 2748
rect 3485 2746 3541 2748
rect 3565 2746 3621 2748
rect 3645 2746 3701 2748
rect 3405 2694 3451 2746
rect 3451 2694 3461 2746
rect 3485 2694 3515 2746
rect 3515 2694 3527 2746
rect 3527 2694 3541 2746
rect 3565 2694 3579 2746
rect 3579 2694 3591 2746
rect 3591 2694 3621 2746
rect 3645 2694 3655 2746
rect 3655 2694 3701 2746
rect 3405 2692 3461 2694
rect 3485 2692 3541 2694
rect 3565 2692 3621 2694
rect 3645 2692 3701 2694
rect 5854 18522 5910 18524
rect 5934 18522 5990 18524
rect 6014 18522 6070 18524
rect 6094 18522 6150 18524
rect 5854 18470 5900 18522
rect 5900 18470 5910 18522
rect 5934 18470 5964 18522
rect 5964 18470 5976 18522
rect 5976 18470 5990 18522
rect 6014 18470 6028 18522
rect 6028 18470 6040 18522
rect 6040 18470 6070 18522
rect 6094 18470 6104 18522
rect 6104 18470 6150 18522
rect 5854 18468 5910 18470
rect 5934 18468 5990 18470
rect 6014 18468 6070 18470
rect 6094 18468 6150 18470
rect 5854 17434 5910 17436
rect 5934 17434 5990 17436
rect 6014 17434 6070 17436
rect 6094 17434 6150 17436
rect 5854 17382 5900 17434
rect 5900 17382 5910 17434
rect 5934 17382 5964 17434
rect 5964 17382 5976 17434
rect 5976 17382 5990 17434
rect 6014 17382 6028 17434
rect 6028 17382 6040 17434
rect 6040 17382 6070 17434
rect 6094 17382 6104 17434
rect 6104 17382 6150 17434
rect 5854 17380 5910 17382
rect 5934 17380 5990 17382
rect 6014 17380 6070 17382
rect 6094 17380 6150 17382
rect 5854 16346 5910 16348
rect 5934 16346 5990 16348
rect 6014 16346 6070 16348
rect 6094 16346 6150 16348
rect 5854 16294 5900 16346
rect 5900 16294 5910 16346
rect 5934 16294 5964 16346
rect 5964 16294 5976 16346
rect 5976 16294 5990 16346
rect 6014 16294 6028 16346
rect 6028 16294 6040 16346
rect 6040 16294 6070 16346
rect 6094 16294 6104 16346
rect 6104 16294 6150 16346
rect 5854 16292 5910 16294
rect 5934 16292 5990 16294
rect 6014 16292 6070 16294
rect 6094 16292 6150 16294
rect 5854 15258 5910 15260
rect 5934 15258 5990 15260
rect 6014 15258 6070 15260
rect 6094 15258 6150 15260
rect 5854 15206 5900 15258
rect 5900 15206 5910 15258
rect 5934 15206 5964 15258
rect 5964 15206 5976 15258
rect 5976 15206 5990 15258
rect 6014 15206 6028 15258
rect 6028 15206 6040 15258
rect 6040 15206 6070 15258
rect 6094 15206 6104 15258
rect 6104 15206 6150 15258
rect 5854 15204 5910 15206
rect 5934 15204 5990 15206
rect 6014 15204 6070 15206
rect 6094 15204 6150 15206
rect 5854 14170 5910 14172
rect 5934 14170 5990 14172
rect 6014 14170 6070 14172
rect 6094 14170 6150 14172
rect 5854 14118 5900 14170
rect 5900 14118 5910 14170
rect 5934 14118 5964 14170
rect 5964 14118 5976 14170
rect 5976 14118 5990 14170
rect 6014 14118 6028 14170
rect 6028 14118 6040 14170
rect 6040 14118 6070 14170
rect 6094 14118 6104 14170
rect 6104 14118 6150 14170
rect 5854 14116 5910 14118
rect 5934 14116 5990 14118
rect 6014 14116 6070 14118
rect 6094 14116 6150 14118
rect 5854 13082 5910 13084
rect 5934 13082 5990 13084
rect 6014 13082 6070 13084
rect 6094 13082 6150 13084
rect 5854 13030 5900 13082
rect 5900 13030 5910 13082
rect 5934 13030 5964 13082
rect 5964 13030 5976 13082
rect 5976 13030 5990 13082
rect 6014 13030 6028 13082
rect 6028 13030 6040 13082
rect 6040 13030 6070 13082
rect 6094 13030 6104 13082
rect 6104 13030 6150 13082
rect 5854 13028 5910 13030
rect 5934 13028 5990 13030
rect 6014 13028 6070 13030
rect 6094 13028 6150 13030
rect 5854 11994 5910 11996
rect 5934 11994 5990 11996
rect 6014 11994 6070 11996
rect 6094 11994 6150 11996
rect 5854 11942 5900 11994
rect 5900 11942 5910 11994
rect 5934 11942 5964 11994
rect 5964 11942 5976 11994
rect 5976 11942 5990 11994
rect 6014 11942 6028 11994
rect 6028 11942 6040 11994
rect 6040 11942 6070 11994
rect 6094 11942 6104 11994
rect 6104 11942 6150 11994
rect 5854 11940 5910 11942
rect 5934 11940 5990 11942
rect 6014 11940 6070 11942
rect 6094 11940 6150 11942
rect 5854 10906 5910 10908
rect 5934 10906 5990 10908
rect 6014 10906 6070 10908
rect 6094 10906 6150 10908
rect 5854 10854 5900 10906
rect 5900 10854 5910 10906
rect 5934 10854 5964 10906
rect 5964 10854 5976 10906
rect 5976 10854 5990 10906
rect 6014 10854 6028 10906
rect 6028 10854 6040 10906
rect 6040 10854 6070 10906
rect 6094 10854 6104 10906
rect 6104 10854 6150 10906
rect 5854 10852 5910 10854
rect 5934 10852 5990 10854
rect 6014 10852 6070 10854
rect 6094 10852 6150 10854
rect 5854 9818 5910 9820
rect 5934 9818 5990 9820
rect 6014 9818 6070 9820
rect 6094 9818 6150 9820
rect 5854 9766 5900 9818
rect 5900 9766 5910 9818
rect 5934 9766 5964 9818
rect 5964 9766 5976 9818
rect 5976 9766 5990 9818
rect 6014 9766 6028 9818
rect 6028 9766 6040 9818
rect 6040 9766 6070 9818
rect 6094 9766 6104 9818
rect 6104 9766 6150 9818
rect 5854 9764 5910 9766
rect 5934 9764 5990 9766
rect 6014 9764 6070 9766
rect 6094 9764 6150 9766
rect 5854 8730 5910 8732
rect 5934 8730 5990 8732
rect 6014 8730 6070 8732
rect 6094 8730 6150 8732
rect 5854 8678 5900 8730
rect 5900 8678 5910 8730
rect 5934 8678 5964 8730
rect 5964 8678 5976 8730
rect 5976 8678 5990 8730
rect 6014 8678 6028 8730
rect 6028 8678 6040 8730
rect 6040 8678 6070 8730
rect 6094 8678 6104 8730
rect 6104 8678 6150 8730
rect 5854 8676 5910 8678
rect 5934 8676 5990 8678
rect 6014 8676 6070 8678
rect 6094 8676 6150 8678
rect 5854 7642 5910 7644
rect 5934 7642 5990 7644
rect 6014 7642 6070 7644
rect 6094 7642 6150 7644
rect 5854 7590 5900 7642
rect 5900 7590 5910 7642
rect 5934 7590 5964 7642
rect 5964 7590 5976 7642
rect 5976 7590 5990 7642
rect 6014 7590 6028 7642
rect 6028 7590 6040 7642
rect 6040 7590 6070 7642
rect 6094 7590 6104 7642
rect 6104 7590 6150 7642
rect 5854 7588 5910 7590
rect 5934 7588 5990 7590
rect 6014 7588 6070 7590
rect 6094 7588 6150 7590
rect 5854 6554 5910 6556
rect 5934 6554 5990 6556
rect 6014 6554 6070 6556
rect 6094 6554 6150 6556
rect 5854 6502 5900 6554
rect 5900 6502 5910 6554
rect 5934 6502 5964 6554
rect 5964 6502 5976 6554
rect 5976 6502 5990 6554
rect 6014 6502 6028 6554
rect 6028 6502 6040 6554
rect 6040 6502 6070 6554
rect 6094 6502 6104 6554
rect 6104 6502 6150 6554
rect 5854 6500 5910 6502
rect 5934 6500 5990 6502
rect 6014 6500 6070 6502
rect 6094 6500 6150 6502
rect 5854 5466 5910 5468
rect 5934 5466 5990 5468
rect 6014 5466 6070 5468
rect 6094 5466 6150 5468
rect 5854 5414 5900 5466
rect 5900 5414 5910 5466
rect 5934 5414 5964 5466
rect 5964 5414 5976 5466
rect 5976 5414 5990 5466
rect 6014 5414 6028 5466
rect 6028 5414 6040 5466
rect 6040 5414 6070 5466
rect 6094 5414 6104 5466
rect 6104 5414 6150 5466
rect 5854 5412 5910 5414
rect 5934 5412 5990 5414
rect 6014 5412 6070 5414
rect 6094 5412 6150 5414
rect 5854 4378 5910 4380
rect 5934 4378 5990 4380
rect 6014 4378 6070 4380
rect 6094 4378 6150 4380
rect 5854 4326 5900 4378
rect 5900 4326 5910 4378
rect 5934 4326 5964 4378
rect 5964 4326 5976 4378
rect 5976 4326 5990 4378
rect 6014 4326 6028 4378
rect 6028 4326 6040 4378
rect 6040 4326 6070 4378
rect 6094 4326 6104 4378
rect 6104 4326 6150 4378
rect 5854 4324 5910 4326
rect 5934 4324 5990 4326
rect 6014 4324 6070 4326
rect 6094 4324 6150 4326
rect 8304 21242 8360 21244
rect 8384 21242 8440 21244
rect 8464 21242 8520 21244
rect 8544 21242 8600 21244
rect 8304 21190 8350 21242
rect 8350 21190 8360 21242
rect 8384 21190 8414 21242
rect 8414 21190 8426 21242
rect 8426 21190 8440 21242
rect 8464 21190 8478 21242
rect 8478 21190 8490 21242
rect 8490 21190 8520 21242
rect 8544 21190 8554 21242
rect 8554 21190 8600 21242
rect 8304 21188 8360 21190
rect 8384 21188 8440 21190
rect 8464 21188 8520 21190
rect 8544 21188 8600 21190
rect 8304 20154 8360 20156
rect 8384 20154 8440 20156
rect 8464 20154 8520 20156
rect 8544 20154 8600 20156
rect 8304 20102 8350 20154
rect 8350 20102 8360 20154
rect 8384 20102 8414 20154
rect 8414 20102 8426 20154
rect 8426 20102 8440 20154
rect 8464 20102 8478 20154
rect 8478 20102 8490 20154
rect 8490 20102 8520 20154
rect 8544 20102 8554 20154
rect 8554 20102 8600 20154
rect 8304 20100 8360 20102
rect 8384 20100 8440 20102
rect 8464 20100 8520 20102
rect 8544 20100 8600 20102
rect 8304 19066 8360 19068
rect 8384 19066 8440 19068
rect 8464 19066 8520 19068
rect 8544 19066 8600 19068
rect 8304 19014 8350 19066
rect 8350 19014 8360 19066
rect 8384 19014 8414 19066
rect 8414 19014 8426 19066
rect 8426 19014 8440 19066
rect 8464 19014 8478 19066
rect 8478 19014 8490 19066
rect 8490 19014 8520 19066
rect 8544 19014 8554 19066
rect 8554 19014 8600 19066
rect 8304 19012 8360 19014
rect 8384 19012 8440 19014
rect 8464 19012 8520 19014
rect 8544 19012 8600 19014
rect 8304 17978 8360 17980
rect 8384 17978 8440 17980
rect 8464 17978 8520 17980
rect 8544 17978 8600 17980
rect 8304 17926 8350 17978
rect 8350 17926 8360 17978
rect 8384 17926 8414 17978
rect 8414 17926 8426 17978
rect 8426 17926 8440 17978
rect 8464 17926 8478 17978
rect 8478 17926 8490 17978
rect 8490 17926 8520 17978
rect 8544 17926 8554 17978
rect 8554 17926 8600 17978
rect 8304 17924 8360 17926
rect 8384 17924 8440 17926
rect 8464 17924 8520 17926
rect 8544 17924 8600 17926
rect 8304 16890 8360 16892
rect 8384 16890 8440 16892
rect 8464 16890 8520 16892
rect 8544 16890 8600 16892
rect 8304 16838 8350 16890
rect 8350 16838 8360 16890
rect 8384 16838 8414 16890
rect 8414 16838 8426 16890
rect 8426 16838 8440 16890
rect 8464 16838 8478 16890
rect 8478 16838 8490 16890
rect 8490 16838 8520 16890
rect 8544 16838 8554 16890
rect 8554 16838 8600 16890
rect 8304 16836 8360 16838
rect 8384 16836 8440 16838
rect 8464 16836 8520 16838
rect 8544 16836 8600 16838
rect 8304 15802 8360 15804
rect 8384 15802 8440 15804
rect 8464 15802 8520 15804
rect 8544 15802 8600 15804
rect 8304 15750 8350 15802
rect 8350 15750 8360 15802
rect 8384 15750 8414 15802
rect 8414 15750 8426 15802
rect 8426 15750 8440 15802
rect 8464 15750 8478 15802
rect 8478 15750 8490 15802
rect 8490 15750 8520 15802
rect 8544 15750 8554 15802
rect 8554 15750 8600 15802
rect 8304 15748 8360 15750
rect 8384 15748 8440 15750
rect 8464 15748 8520 15750
rect 8544 15748 8600 15750
rect 8304 14714 8360 14716
rect 8384 14714 8440 14716
rect 8464 14714 8520 14716
rect 8544 14714 8600 14716
rect 8304 14662 8350 14714
rect 8350 14662 8360 14714
rect 8384 14662 8414 14714
rect 8414 14662 8426 14714
rect 8426 14662 8440 14714
rect 8464 14662 8478 14714
rect 8478 14662 8490 14714
rect 8490 14662 8520 14714
rect 8544 14662 8554 14714
rect 8554 14662 8600 14714
rect 8304 14660 8360 14662
rect 8384 14660 8440 14662
rect 8464 14660 8520 14662
rect 8544 14660 8600 14662
rect 8304 13626 8360 13628
rect 8384 13626 8440 13628
rect 8464 13626 8520 13628
rect 8544 13626 8600 13628
rect 8304 13574 8350 13626
rect 8350 13574 8360 13626
rect 8384 13574 8414 13626
rect 8414 13574 8426 13626
rect 8426 13574 8440 13626
rect 8464 13574 8478 13626
rect 8478 13574 8490 13626
rect 8490 13574 8520 13626
rect 8544 13574 8554 13626
rect 8554 13574 8600 13626
rect 8304 13572 8360 13574
rect 8384 13572 8440 13574
rect 8464 13572 8520 13574
rect 8544 13572 8600 13574
rect 8304 12538 8360 12540
rect 8384 12538 8440 12540
rect 8464 12538 8520 12540
rect 8544 12538 8600 12540
rect 8304 12486 8350 12538
rect 8350 12486 8360 12538
rect 8384 12486 8414 12538
rect 8414 12486 8426 12538
rect 8426 12486 8440 12538
rect 8464 12486 8478 12538
rect 8478 12486 8490 12538
rect 8490 12486 8520 12538
rect 8544 12486 8554 12538
rect 8554 12486 8600 12538
rect 8304 12484 8360 12486
rect 8384 12484 8440 12486
rect 8464 12484 8520 12486
rect 8544 12484 8600 12486
rect 8304 11450 8360 11452
rect 8384 11450 8440 11452
rect 8464 11450 8520 11452
rect 8544 11450 8600 11452
rect 8304 11398 8350 11450
rect 8350 11398 8360 11450
rect 8384 11398 8414 11450
rect 8414 11398 8426 11450
rect 8426 11398 8440 11450
rect 8464 11398 8478 11450
rect 8478 11398 8490 11450
rect 8490 11398 8520 11450
rect 8544 11398 8554 11450
rect 8554 11398 8600 11450
rect 8304 11396 8360 11398
rect 8384 11396 8440 11398
rect 8464 11396 8520 11398
rect 8544 11396 8600 11398
rect 8304 10362 8360 10364
rect 8384 10362 8440 10364
rect 8464 10362 8520 10364
rect 8544 10362 8600 10364
rect 8304 10310 8350 10362
rect 8350 10310 8360 10362
rect 8384 10310 8414 10362
rect 8414 10310 8426 10362
rect 8426 10310 8440 10362
rect 8464 10310 8478 10362
rect 8478 10310 8490 10362
rect 8490 10310 8520 10362
rect 8544 10310 8554 10362
rect 8554 10310 8600 10362
rect 8304 10308 8360 10310
rect 8384 10308 8440 10310
rect 8464 10308 8520 10310
rect 8544 10308 8600 10310
rect 8304 9274 8360 9276
rect 8384 9274 8440 9276
rect 8464 9274 8520 9276
rect 8544 9274 8600 9276
rect 8304 9222 8350 9274
rect 8350 9222 8360 9274
rect 8384 9222 8414 9274
rect 8414 9222 8426 9274
rect 8426 9222 8440 9274
rect 8464 9222 8478 9274
rect 8478 9222 8490 9274
rect 8490 9222 8520 9274
rect 8544 9222 8554 9274
rect 8554 9222 8600 9274
rect 8304 9220 8360 9222
rect 8384 9220 8440 9222
rect 8464 9220 8520 9222
rect 8544 9220 8600 9222
rect 8304 8186 8360 8188
rect 8384 8186 8440 8188
rect 8464 8186 8520 8188
rect 8544 8186 8600 8188
rect 8304 8134 8350 8186
rect 8350 8134 8360 8186
rect 8384 8134 8414 8186
rect 8414 8134 8426 8186
rect 8426 8134 8440 8186
rect 8464 8134 8478 8186
rect 8478 8134 8490 8186
rect 8490 8134 8520 8186
rect 8544 8134 8554 8186
rect 8554 8134 8600 8186
rect 8304 8132 8360 8134
rect 8384 8132 8440 8134
rect 8464 8132 8520 8134
rect 8544 8132 8600 8134
rect 8304 7098 8360 7100
rect 8384 7098 8440 7100
rect 8464 7098 8520 7100
rect 8544 7098 8600 7100
rect 8304 7046 8350 7098
rect 8350 7046 8360 7098
rect 8384 7046 8414 7098
rect 8414 7046 8426 7098
rect 8426 7046 8440 7098
rect 8464 7046 8478 7098
rect 8478 7046 8490 7098
rect 8490 7046 8520 7098
rect 8544 7046 8554 7098
rect 8554 7046 8600 7098
rect 8304 7044 8360 7046
rect 8384 7044 8440 7046
rect 8464 7044 8520 7046
rect 8544 7044 8600 7046
rect 8304 6010 8360 6012
rect 8384 6010 8440 6012
rect 8464 6010 8520 6012
rect 8544 6010 8600 6012
rect 8304 5958 8350 6010
rect 8350 5958 8360 6010
rect 8384 5958 8414 6010
rect 8414 5958 8426 6010
rect 8426 5958 8440 6010
rect 8464 5958 8478 6010
rect 8478 5958 8490 6010
rect 8490 5958 8520 6010
rect 8544 5958 8554 6010
rect 8554 5958 8600 6010
rect 8304 5956 8360 5958
rect 8384 5956 8440 5958
rect 8464 5956 8520 5958
rect 8544 5956 8600 5958
rect 8304 4922 8360 4924
rect 8384 4922 8440 4924
rect 8464 4922 8520 4924
rect 8544 4922 8600 4924
rect 8304 4870 8350 4922
rect 8350 4870 8360 4922
rect 8384 4870 8414 4922
rect 8414 4870 8426 4922
rect 8426 4870 8440 4922
rect 8464 4870 8478 4922
rect 8478 4870 8490 4922
rect 8490 4870 8520 4922
rect 8544 4870 8554 4922
rect 8554 4870 8600 4922
rect 8304 4868 8360 4870
rect 8384 4868 8440 4870
rect 8464 4868 8520 4870
rect 8544 4868 8600 4870
rect 5854 3290 5910 3292
rect 5934 3290 5990 3292
rect 6014 3290 6070 3292
rect 6094 3290 6150 3292
rect 5854 3238 5900 3290
rect 5900 3238 5910 3290
rect 5934 3238 5964 3290
rect 5964 3238 5976 3290
rect 5976 3238 5990 3290
rect 6014 3238 6028 3290
rect 6028 3238 6040 3290
rect 6040 3238 6070 3290
rect 6094 3238 6104 3290
rect 6104 3238 6150 3290
rect 5854 3236 5910 3238
rect 5934 3236 5990 3238
rect 6014 3236 6070 3238
rect 6094 3236 6150 3238
rect 8304 3834 8360 3836
rect 8384 3834 8440 3836
rect 8464 3834 8520 3836
rect 8544 3834 8600 3836
rect 8304 3782 8350 3834
rect 8350 3782 8360 3834
rect 8384 3782 8414 3834
rect 8414 3782 8426 3834
rect 8426 3782 8440 3834
rect 8464 3782 8478 3834
rect 8478 3782 8490 3834
rect 8490 3782 8520 3834
rect 8544 3782 8554 3834
rect 8554 3782 8600 3834
rect 8304 3780 8360 3782
rect 8384 3780 8440 3782
rect 8464 3780 8520 3782
rect 8544 3780 8600 3782
rect 8304 2746 8360 2748
rect 8384 2746 8440 2748
rect 8464 2746 8520 2748
rect 8544 2746 8600 2748
rect 8304 2694 8350 2746
rect 8350 2694 8360 2746
rect 8384 2694 8414 2746
rect 8414 2694 8426 2746
rect 8426 2694 8440 2746
rect 8464 2694 8478 2746
rect 8478 2694 8490 2746
rect 8490 2694 8520 2746
rect 8544 2694 8554 2746
rect 8554 2694 8600 2746
rect 8304 2692 8360 2694
rect 8384 2692 8440 2694
rect 8464 2692 8520 2694
rect 8544 2692 8600 2694
rect 10753 20698 10809 20700
rect 10833 20698 10889 20700
rect 10913 20698 10969 20700
rect 10993 20698 11049 20700
rect 10753 20646 10799 20698
rect 10799 20646 10809 20698
rect 10833 20646 10863 20698
rect 10863 20646 10875 20698
rect 10875 20646 10889 20698
rect 10913 20646 10927 20698
rect 10927 20646 10939 20698
rect 10939 20646 10969 20698
rect 10993 20646 11003 20698
rect 11003 20646 11049 20698
rect 10753 20644 10809 20646
rect 10833 20644 10889 20646
rect 10913 20644 10969 20646
rect 10993 20644 11049 20646
rect 10753 19610 10809 19612
rect 10833 19610 10889 19612
rect 10913 19610 10969 19612
rect 10993 19610 11049 19612
rect 10753 19558 10799 19610
rect 10799 19558 10809 19610
rect 10833 19558 10863 19610
rect 10863 19558 10875 19610
rect 10875 19558 10889 19610
rect 10913 19558 10927 19610
rect 10927 19558 10939 19610
rect 10939 19558 10969 19610
rect 10993 19558 11003 19610
rect 11003 19558 11049 19610
rect 10753 19556 10809 19558
rect 10833 19556 10889 19558
rect 10913 19556 10969 19558
rect 10993 19556 11049 19558
rect 10753 18522 10809 18524
rect 10833 18522 10889 18524
rect 10913 18522 10969 18524
rect 10993 18522 11049 18524
rect 10753 18470 10799 18522
rect 10799 18470 10809 18522
rect 10833 18470 10863 18522
rect 10863 18470 10875 18522
rect 10875 18470 10889 18522
rect 10913 18470 10927 18522
rect 10927 18470 10939 18522
rect 10939 18470 10969 18522
rect 10993 18470 11003 18522
rect 11003 18470 11049 18522
rect 10753 18468 10809 18470
rect 10833 18468 10889 18470
rect 10913 18468 10969 18470
rect 10993 18468 11049 18470
rect 13203 21242 13259 21244
rect 13283 21242 13339 21244
rect 13363 21242 13419 21244
rect 13443 21242 13499 21244
rect 13203 21190 13249 21242
rect 13249 21190 13259 21242
rect 13283 21190 13313 21242
rect 13313 21190 13325 21242
rect 13325 21190 13339 21242
rect 13363 21190 13377 21242
rect 13377 21190 13389 21242
rect 13389 21190 13419 21242
rect 13443 21190 13453 21242
rect 13453 21190 13499 21242
rect 13203 21188 13259 21190
rect 13283 21188 13339 21190
rect 13363 21188 13419 21190
rect 13443 21188 13499 21190
rect 13203 20154 13259 20156
rect 13283 20154 13339 20156
rect 13363 20154 13419 20156
rect 13443 20154 13499 20156
rect 13203 20102 13249 20154
rect 13249 20102 13259 20154
rect 13283 20102 13313 20154
rect 13313 20102 13325 20154
rect 13325 20102 13339 20154
rect 13363 20102 13377 20154
rect 13377 20102 13389 20154
rect 13389 20102 13419 20154
rect 13443 20102 13453 20154
rect 13453 20102 13499 20154
rect 13203 20100 13259 20102
rect 13283 20100 13339 20102
rect 13363 20100 13419 20102
rect 13443 20100 13499 20102
rect 13203 19066 13259 19068
rect 13283 19066 13339 19068
rect 13363 19066 13419 19068
rect 13443 19066 13499 19068
rect 13203 19014 13249 19066
rect 13249 19014 13259 19066
rect 13283 19014 13313 19066
rect 13313 19014 13325 19066
rect 13325 19014 13339 19066
rect 13363 19014 13377 19066
rect 13377 19014 13389 19066
rect 13389 19014 13419 19066
rect 13443 19014 13453 19066
rect 13453 19014 13499 19066
rect 13203 19012 13259 19014
rect 13283 19012 13339 19014
rect 13363 19012 13419 19014
rect 13443 19012 13499 19014
rect 10753 17434 10809 17436
rect 10833 17434 10889 17436
rect 10913 17434 10969 17436
rect 10993 17434 11049 17436
rect 10753 17382 10799 17434
rect 10799 17382 10809 17434
rect 10833 17382 10863 17434
rect 10863 17382 10875 17434
rect 10875 17382 10889 17434
rect 10913 17382 10927 17434
rect 10927 17382 10939 17434
rect 10939 17382 10969 17434
rect 10993 17382 11003 17434
rect 11003 17382 11049 17434
rect 10753 17380 10809 17382
rect 10833 17380 10889 17382
rect 10913 17380 10969 17382
rect 10993 17380 11049 17382
rect 10753 16346 10809 16348
rect 10833 16346 10889 16348
rect 10913 16346 10969 16348
rect 10993 16346 11049 16348
rect 10753 16294 10799 16346
rect 10799 16294 10809 16346
rect 10833 16294 10863 16346
rect 10863 16294 10875 16346
rect 10875 16294 10889 16346
rect 10913 16294 10927 16346
rect 10927 16294 10939 16346
rect 10939 16294 10969 16346
rect 10993 16294 11003 16346
rect 11003 16294 11049 16346
rect 10753 16292 10809 16294
rect 10833 16292 10889 16294
rect 10913 16292 10969 16294
rect 10993 16292 11049 16294
rect 10753 15258 10809 15260
rect 10833 15258 10889 15260
rect 10913 15258 10969 15260
rect 10993 15258 11049 15260
rect 10753 15206 10799 15258
rect 10799 15206 10809 15258
rect 10833 15206 10863 15258
rect 10863 15206 10875 15258
rect 10875 15206 10889 15258
rect 10913 15206 10927 15258
rect 10927 15206 10939 15258
rect 10939 15206 10969 15258
rect 10993 15206 11003 15258
rect 11003 15206 11049 15258
rect 10753 15204 10809 15206
rect 10833 15204 10889 15206
rect 10913 15204 10969 15206
rect 10993 15204 11049 15206
rect 13203 17978 13259 17980
rect 13283 17978 13339 17980
rect 13363 17978 13419 17980
rect 13443 17978 13499 17980
rect 13203 17926 13249 17978
rect 13249 17926 13259 17978
rect 13283 17926 13313 17978
rect 13313 17926 13325 17978
rect 13325 17926 13339 17978
rect 13363 17926 13377 17978
rect 13377 17926 13389 17978
rect 13389 17926 13419 17978
rect 13443 17926 13453 17978
rect 13453 17926 13499 17978
rect 13203 17924 13259 17926
rect 13283 17924 13339 17926
rect 13363 17924 13419 17926
rect 13443 17924 13499 17926
rect 13203 16890 13259 16892
rect 13283 16890 13339 16892
rect 13363 16890 13419 16892
rect 13443 16890 13499 16892
rect 13203 16838 13249 16890
rect 13249 16838 13259 16890
rect 13283 16838 13313 16890
rect 13313 16838 13325 16890
rect 13325 16838 13339 16890
rect 13363 16838 13377 16890
rect 13377 16838 13389 16890
rect 13389 16838 13419 16890
rect 13443 16838 13453 16890
rect 13453 16838 13499 16890
rect 13203 16836 13259 16838
rect 13283 16836 13339 16838
rect 13363 16836 13419 16838
rect 13443 16836 13499 16838
rect 13203 15802 13259 15804
rect 13283 15802 13339 15804
rect 13363 15802 13419 15804
rect 13443 15802 13499 15804
rect 13203 15750 13249 15802
rect 13249 15750 13259 15802
rect 13283 15750 13313 15802
rect 13313 15750 13325 15802
rect 13325 15750 13339 15802
rect 13363 15750 13377 15802
rect 13377 15750 13389 15802
rect 13389 15750 13419 15802
rect 13443 15750 13453 15802
rect 13453 15750 13499 15802
rect 13203 15748 13259 15750
rect 13283 15748 13339 15750
rect 13363 15748 13419 15750
rect 13443 15748 13499 15750
rect 13203 14714 13259 14716
rect 13283 14714 13339 14716
rect 13363 14714 13419 14716
rect 13443 14714 13499 14716
rect 13203 14662 13249 14714
rect 13249 14662 13259 14714
rect 13283 14662 13313 14714
rect 13313 14662 13325 14714
rect 13325 14662 13339 14714
rect 13363 14662 13377 14714
rect 13377 14662 13389 14714
rect 13389 14662 13419 14714
rect 13443 14662 13453 14714
rect 13453 14662 13499 14714
rect 13203 14660 13259 14662
rect 13283 14660 13339 14662
rect 13363 14660 13419 14662
rect 13443 14660 13499 14662
rect 10753 14170 10809 14172
rect 10833 14170 10889 14172
rect 10913 14170 10969 14172
rect 10993 14170 11049 14172
rect 10753 14118 10799 14170
rect 10799 14118 10809 14170
rect 10833 14118 10863 14170
rect 10863 14118 10875 14170
rect 10875 14118 10889 14170
rect 10913 14118 10927 14170
rect 10927 14118 10939 14170
rect 10939 14118 10969 14170
rect 10993 14118 11003 14170
rect 11003 14118 11049 14170
rect 10753 14116 10809 14118
rect 10833 14116 10889 14118
rect 10913 14116 10969 14118
rect 10993 14116 11049 14118
rect 10753 13082 10809 13084
rect 10833 13082 10889 13084
rect 10913 13082 10969 13084
rect 10993 13082 11049 13084
rect 10753 13030 10799 13082
rect 10799 13030 10809 13082
rect 10833 13030 10863 13082
rect 10863 13030 10875 13082
rect 10875 13030 10889 13082
rect 10913 13030 10927 13082
rect 10927 13030 10939 13082
rect 10939 13030 10969 13082
rect 10993 13030 11003 13082
rect 11003 13030 11049 13082
rect 10753 13028 10809 13030
rect 10833 13028 10889 13030
rect 10913 13028 10969 13030
rect 10993 13028 11049 13030
rect 10753 11994 10809 11996
rect 10833 11994 10889 11996
rect 10913 11994 10969 11996
rect 10993 11994 11049 11996
rect 10753 11942 10799 11994
rect 10799 11942 10809 11994
rect 10833 11942 10863 11994
rect 10863 11942 10875 11994
rect 10875 11942 10889 11994
rect 10913 11942 10927 11994
rect 10927 11942 10939 11994
rect 10939 11942 10969 11994
rect 10993 11942 11003 11994
rect 11003 11942 11049 11994
rect 10753 11940 10809 11942
rect 10833 11940 10889 11942
rect 10913 11940 10969 11942
rect 10993 11940 11049 11942
rect 10753 10906 10809 10908
rect 10833 10906 10889 10908
rect 10913 10906 10969 10908
rect 10993 10906 11049 10908
rect 10753 10854 10799 10906
rect 10799 10854 10809 10906
rect 10833 10854 10863 10906
rect 10863 10854 10875 10906
rect 10875 10854 10889 10906
rect 10913 10854 10927 10906
rect 10927 10854 10939 10906
rect 10939 10854 10969 10906
rect 10993 10854 11003 10906
rect 11003 10854 11049 10906
rect 10753 10852 10809 10854
rect 10833 10852 10889 10854
rect 10913 10852 10969 10854
rect 10993 10852 11049 10854
rect 10753 9818 10809 9820
rect 10833 9818 10889 9820
rect 10913 9818 10969 9820
rect 10993 9818 11049 9820
rect 10753 9766 10799 9818
rect 10799 9766 10809 9818
rect 10833 9766 10863 9818
rect 10863 9766 10875 9818
rect 10875 9766 10889 9818
rect 10913 9766 10927 9818
rect 10927 9766 10939 9818
rect 10939 9766 10969 9818
rect 10993 9766 11003 9818
rect 11003 9766 11049 9818
rect 10753 9764 10809 9766
rect 10833 9764 10889 9766
rect 10913 9764 10969 9766
rect 10993 9764 11049 9766
rect 10753 8730 10809 8732
rect 10833 8730 10889 8732
rect 10913 8730 10969 8732
rect 10993 8730 11049 8732
rect 10753 8678 10799 8730
rect 10799 8678 10809 8730
rect 10833 8678 10863 8730
rect 10863 8678 10875 8730
rect 10875 8678 10889 8730
rect 10913 8678 10927 8730
rect 10927 8678 10939 8730
rect 10939 8678 10969 8730
rect 10993 8678 11003 8730
rect 11003 8678 11049 8730
rect 10753 8676 10809 8678
rect 10833 8676 10889 8678
rect 10913 8676 10969 8678
rect 10993 8676 11049 8678
rect 10753 7642 10809 7644
rect 10833 7642 10889 7644
rect 10913 7642 10969 7644
rect 10993 7642 11049 7644
rect 10753 7590 10799 7642
rect 10799 7590 10809 7642
rect 10833 7590 10863 7642
rect 10863 7590 10875 7642
rect 10875 7590 10889 7642
rect 10913 7590 10927 7642
rect 10927 7590 10939 7642
rect 10939 7590 10969 7642
rect 10993 7590 11003 7642
rect 11003 7590 11049 7642
rect 10753 7588 10809 7590
rect 10833 7588 10889 7590
rect 10913 7588 10969 7590
rect 10993 7588 11049 7590
rect 10753 6554 10809 6556
rect 10833 6554 10889 6556
rect 10913 6554 10969 6556
rect 10993 6554 11049 6556
rect 10753 6502 10799 6554
rect 10799 6502 10809 6554
rect 10833 6502 10863 6554
rect 10863 6502 10875 6554
rect 10875 6502 10889 6554
rect 10913 6502 10927 6554
rect 10927 6502 10939 6554
rect 10939 6502 10969 6554
rect 10993 6502 11003 6554
rect 11003 6502 11049 6554
rect 10753 6500 10809 6502
rect 10833 6500 10889 6502
rect 10913 6500 10969 6502
rect 10993 6500 11049 6502
rect 10753 5466 10809 5468
rect 10833 5466 10889 5468
rect 10913 5466 10969 5468
rect 10993 5466 11049 5468
rect 10753 5414 10799 5466
rect 10799 5414 10809 5466
rect 10833 5414 10863 5466
rect 10863 5414 10875 5466
rect 10875 5414 10889 5466
rect 10913 5414 10927 5466
rect 10927 5414 10939 5466
rect 10939 5414 10969 5466
rect 10993 5414 11003 5466
rect 11003 5414 11049 5466
rect 10753 5412 10809 5414
rect 10833 5412 10889 5414
rect 10913 5412 10969 5414
rect 10993 5412 11049 5414
rect 10753 4378 10809 4380
rect 10833 4378 10889 4380
rect 10913 4378 10969 4380
rect 10993 4378 11049 4380
rect 10753 4326 10799 4378
rect 10799 4326 10809 4378
rect 10833 4326 10863 4378
rect 10863 4326 10875 4378
rect 10875 4326 10889 4378
rect 10913 4326 10927 4378
rect 10927 4326 10939 4378
rect 10939 4326 10969 4378
rect 10993 4326 11003 4378
rect 11003 4326 11049 4378
rect 10753 4324 10809 4326
rect 10833 4324 10889 4326
rect 10913 4324 10969 4326
rect 10993 4324 11049 4326
rect 13203 13626 13259 13628
rect 13283 13626 13339 13628
rect 13363 13626 13419 13628
rect 13443 13626 13499 13628
rect 13203 13574 13249 13626
rect 13249 13574 13259 13626
rect 13283 13574 13313 13626
rect 13313 13574 13325 13626
rect 13325 13574 13339 13626
rect 13363 13574 13377 13626
rect 13377 13574 13389 13626
rect 13389 13574 13419 13626
rect 13443 13574 13453 13626
rect 13453 13574 13499 13626
rect 13203 13572 13259 13574
rect 13283 13572 13339 13574
rect 13363 13572 13419 13574
rect 13443 13572 13499 13574
rect 13203 12538 13259 12540
rect 13283 12538 13339 12540
rect 13363 12538 13419 12540
rect 13443 12538 13499 12540
rect 13203 12486 13249 12538
rect 13249 12486 13259 12538
rect 13283 12486 13313 12538
rect 13313 12486 13325 12538
rect 13325 12486 13339 12538
rect 13363 12486 13377 12538
rect 13377 12486 13389 12538
rect 13389 12486 13419 12538
rect 13443 12486 13453 12538
rect 13453 12486 13499 12538
rect 13203 12484 13259 12486
rect 13283 12484 13339 12486
rect 13363 12484 13419 12486
rect 13443 12484 13499 12486
rect 13203 11450 13259 11452
rect 13283 11450 13339 11452
rect 13363 11450 13419 11452
rect 13443 11450 13499 11452
rect 13203 11398 13249 11450
rect 13249 11398 13259 11450
rect 13283 11398 13313 11450
rect 13313 11398 13325 11450
rect 13325 11398 13339 11450
rect 13363 11398 13377 11450
rect 13377 11398 13389 11450
rect 13389 11398 13419 11450
rect 13443 11398 13453 11450
rect 13453 11398 13499 11450
rect 13203 11396 13259 11398
rect 13283 11396 13339 11398
rect 13363 11396 13419 11398
rect 13443 11396 13499 11398
rect 15652 20698 15708 20700
rect 15732 20698 15788 20700
rect 15812 20698 15868 20700
rect 15892 20698 15948 20700
rect 15652 20646 15698 20698
rect 15698 20646 15708 20698
rect 15732 20646 15762 20698
rect 15762 20646 15774 20698
rect 15774 20646 15788 20698
rect 15812 20646 15826 20698
rect 15826 20646 15838 20698
rect 15838 20646 15868 20698
rect 15892 20646 15902 20698
rect 15902 20646 15948 20698
rect 15652 20644 15708 20646
rect 15732 20644 15788 20646
rect 15812 20644 15868 20646
rect 15892 20644 15948 20646
rect 15652 19610 15708 19612
rect 15732 19610 15788 19612
rect 15812 19610 15868 19612
rect 15892 19610 15948 19612
rect 15652 19558 15698 19610
rect 15698 19558 15708 19610
rect 15732 19558 15762 19610
rect 15762 19558 15774 19610
rect 15774 19558 15788 19610
rect 15812 19558 15826 19610
rect 15826 19558 15838 19610
rect 15838 19558 15868 19610
rect 15892 19558 15902 19610
rect 15902 19558 15948 19610
rect 15652 19556 15708 19558
rect 15732 19556 15788 19558
rect 15812 19556 15868 19558
rect 15892 19556 15948 19558
rect 15652 18522 15708 18524
rect 15732 18522 15788 18524
rect 15812 18522 15868 18524
rect 15892 18522 15948 18524
rect 15652 18470 15698 18522
rect 15698 18470 15708 18522
rect 15732 18470 15762 18522
rect 15762 18470 15774 18522
rect 15774 18470 15788 18522
rect 15812 18470 15826 18522
rect 15826 18470 15838 18522
rect 15838 18470 15868 18522
rect 15892 18470 15902 18522
rect 15902 18470 15948 18522
rect 15652 18468 15708 18470
rect 15732 18468 15788 18470
rect 15812 18468 15868 18470
rect 15892 18468 15948 18470
rect 15652 17434 15708 17436
rect 15732 17434 15788 17436
rect 15812 17434 15868 17436
rect 15892 17434 15948 17436
rect 15652 17382 15698 17434
rect 15698 17382 15708 17434
rect 15732 17382 15762 17434
rect 15762 17382 15774 17434
rect 15774 17382 15788 17434
rect 15812 17382 15826 17434
rect 15826 17382 15838 17434
rect 15838 17382 15868 17434
rect 15892 17382 15902 17434
rect 15902 17382 15948 17434
rect 15652 17380 15708 17382
rect 15732 17380 15788 17382
rect 15812 17380 15868 17382
rect 15892 17380 15948 17382
rect 15652 16346 15708 16348
rect 15732 16346 15788 16348
rect 15812 16346 15868 16348
rect 15892 16346 15948 16348
rect 15652 16294 15698 16346
rect 15698 16294 15708 16346
rect 15732 16294 15762 16346
rect 15762 16294 15774 16346
rect 15774 16294 15788 16346
rect 15812 16294 15826 16346
rect 15826 16294 15838 16346
rect 15838 16294 15868 16346
rect 15892 16294 15902 16346
rect 15902 16294 15948 16346
rect 15652 16292 15708 16294
rect 15732 16292 15788 16294
rect 15812 16292 15868 16294
rect 15892 16292 15948 16294
rect 15652 15258 15708 15260
rect 15732 15258 15788 15260
rect 15812 15258 15868 15260
rect 15892 15258 15948 15260
rect 15652 15206 15698 15258
rect 15698 15206 15708 15258
rect 15732 15206 15762 15258
rect 15762 15206 15774 15258
rect 15774 15206 15788 15258
rect 15812 15206 15826 15258
rect 15826 15206 15838 15258
rect 15838 15206 15868 15258
rect 15892 15206 15902 15258
rect 15902 15206 15948 15258
rect 15652 15204 15708 15206
rect 15732 15204 15788 15206
rect 15812 15204 15868 15206
rect 15892 15204 15948 15206
rect 13203 10362 13259 10364
rect 13283 10362 13339 10364
rect 13363 10362 13419 10364
rect 13443 10362 13499 10364
rect 13203 10310 13249 10362
rect 13249 10310 13259 10362
rect 13283 10310 13313 10362
rect 13313 10310 13325 10362
rect 13325 10310 13339 10362
rect 13363 10310 13377 10362
rect 13377 10310 13389 10362
rect 13389 10310 13419 10362
rect 13443 10310 13453 10362
rect 13453 10310 13499 10362
rect 13203 10308 13259 10310
rect 13283 10308 13339 10310
rect 13363 10308 13419 10310
rect 13443 10308 13499 10310
rect 13203 9274 13259 9276
rect 13283 9274 13339 9276
rect 13363 9274 13419 9276
rect 13443 9274 13499 9276
rect 13203 9222 13249 9274
rect 13249 9222 13259 9274
rect 13283 9222 13313 9274
rect 13313 9222 13325 9274
rect 13325 9222 13339 9274
rect 13363 9222 13377 9274
rect 13377 9222 13389 9274
rect 13389 9222 13419 9274
rect 13443 9222 13453 9274
rect 13453 9222 13499 9274
rect 13203 9220 13259 9222
rect 13283 9220 13339 9222
rect 13363 9220 13419 9222
rect 13443 9220 13499 9222
rect 13203 8186 13259 8188
rect 13283 8186 13339 8188
rect 13363 8186 13419 8188
rect 13443 8186 13499 8188
rect 13203 8134 13249 8186
rect 13249 8134 13259 8186
rect 13283 8134 13313 8186
rect 13313 8134 13325 8186
rect 13325 8134 13339 8186
rect 13363 8134 13377 8186
rect 13377 8134 13389 8186
rect 13389 8134 13419 8186
rect 13443 8134 13453 8186
rect 13453 8134 13499 8186
rect 13203 8132 13259 8134
rect 13283 8132 13339 8134
rect 13363 8132 13419 8134
rect 13443 8132 13499 8134
rect 13203 7098 13259 7100
rect 13283 7098 13339 7100
rect 13363 7098 13419 7100
rect 13443 7098 13499 7100
rect 13203 7046 13249 7098
rect 13249 7046 13259 7098
rect 13283 7046 13313 7098
rect 13313 7046 13325 7098
rect 13325 7046 13339 7098
rect 13363 7046 13377 7098
rect 13377 7046 13389 7098
rect 13389 7046 13419 7098
rect 13443 7046 13453 7098
rect 13453 7046 13499 7098
rect 13203 7044 13259 7046
rect 13283 7044 13339 7046
rect 13363 7044 13419 7046
rect 13443 7044 13499 7046
rect 13203 6010 13259 6012
rect 13283 6010 13339 6012
rect 13363 6010 13419 6012
rect 13443 6010 13499 6012
rect 13203 5958 13249 6010
rect 13249 5958 13259 6010
rect 13283 5958 13313 6010
rect 13313 5958 13325 6010
rect 13325 5958 13339 6010
rect 13363 5958 13377 6010
rect 13377 5958 13389 6010
rect 13389 5958 13419 6010
rect 13443 5958 13453 6010
rect 13453 5958 13499 6010
rect 13203 5956 13259 5958
rect 13283 5956 13339 5958
rect 13363 5956 13419 5958
rect 13443 5956 13499 5958
rect 10753 3290 10809 3292
rect 10833 3290 10889 3292
rect 10913 3290 10969 3292
rect 10993 3290 11049 3292
rect 10753 3238 10799 3290
rect 10799 3238 10809 3290
rect 10833 3238 10863 3290
rect 10863 3238 10875 3290
rect 10875 3238 10889 3290
rect 10913 3238 10927 3290
rect 10927 3238 10939 3290
rect 10939 3238 10969 3290
rect 10993 3238 11003 3290
rect 11003 3238 11049 3290
rect 10753 3236 10809 3238
rect 10833 3236 10889 3238
rect 10913 3236 10969 3238
rect 10993 3236 11049 3238
rect 13203 4922 13259 4924
rect 13283 4922 13339 4924
rect 13363 4922 13419 4924
rect 13443 4922 13499 4924
rect 13203 4870 13249 4922
rect 13249 4870 13259 4922
rect 13283 4870 13313 4922
rect 13313 4870 13325 4922
rect 13325 4870 13339 4922
rect 13363 4870 13377 4922
rect 13377 4870 13389 4922
rect 13389 4870 13419 4922
rect 13443 4870 13453 4922
rect 13453 4870 13499 4922
rect 13203 4868 13259 4870
rect 13283 4868 13339 4870
rect 13363 4868 13419 4870
rect 13443 4868 13499 4870
rect 13203 3834 13259 3836
rect 13283 3834 13339 3836
rect 13363 3834 13419 3836
rect 13443 3834 13499 3836
rect 13203 3782 13249 3834
rect 13249 3782 13259 3834
rect 13283 3782 13313 3834
rect 13313 3782 13325 3834
rect 13325 3782 13339 3834
rect 13363 3782 13377 3834
rect 13377 3782 13389 3834
rect 13389 3782 13419 3834
rect 13443 3782 13453 3834
rect 13453 3782 13499 3834
rect 13203 3780 13259 3782
rect 13283 3780 13339 3782
rect 13363 3780 13419 3782
rect 13443 3780 13499 3782
rect 13203 2746 13259 2748
rect 13283 2746 13339 2748
rect 13363 2746 13419 2748
rect 13443 2746 13499 2748
rect 13203 2694 13249 2746
rect 13249 2694 13259 2746
rect 13283 2694 13313 2746
rect 13313 2694 13325 2746
rect 13325 2694 13339 2746
rect 13363 2694 13377 2746
rect 13377 2694 13389 2746
rect 13389 2694 13419 2746
rect 13443 2694 13453 2746
rect 13453 2694 13499 2746
rect 13203 2692 13259 2694
rect 13283 2692 13339 2694
rect 13363 2692 13419 2694
rect 13443 2692 13499 2694
rect 15652 14170 15708 14172
rect 15732 14170 15788 14172
rect 15812 14170 15868 14172
rect 15892 14170 15948 14172
rect 15652 14118 15698 14170
rect 15698 14118 15708 14170
rect 15732 14118 15762 14170
rect 15762 14118 15774 14170
rect 15774 14118 15788 14170
rect 15812 14118 15826 14170
rect 15826 14118 15838 14170
rect 15838 14118 15868 14170
rect 15892 14118 15902 14170
rect 15902 14118 15948 14170
rect 15652 14116 15708 14118
rect 15732 14116 15788 14118
rect 15812 14116 15868 14118
rect 15892 14116 15948 14118
rect 18102 21242 18158 21244
rect 18182 21242 18238 21244
rect 18262 21242 18318 21244
rect 18342 21242 18398 21244
rect 18102 21190 18148 21242
rect 18148 21190 18158 21242
rect 18182 21190 18212 21242
rect 18212 21190 18224 21242
rect 18224 21190 18238 21242
rect 18262 21190 18276 21242
rect 18276 21190 18288 21242
rect 18288 21190 18318 21242
rect 18342 21190 18352 21242
rect 18352 21190 18398 21242
rect 18102 21188 18158 21190
rect 18182 21188 18238 21190
rect 18262 21188 18318 21190
rect 18342 21188 18398 21190
rect 18102 20154 18158 20156
rect 18182 20154 18238 20156
rect 18262 20154 18318 20156
rect 18342 20154 18398 20156
rect 18102 20102 18148 20154
rect 18148 20102 18158 20154
rect 18182 20102 18212 20154
rect 18212 20102 18224 20154
rect 18224 20102 18238 20154
rect 18262 20102 18276 20154
rect 18276 20102 18288 20154
rect 18288 20102 18318 20154
rect 18342 20102 18352 20154
rect 18352 20102 18398 20154
rect 18102 20100 18158 20102
rect 18182 20100 18238 20102
rect 18262 20100 18318 20102
rect 18342 20100 18398 20102
rect 20551 21786 20607 21788
rect 20631 21786 20687 21788
rect 20711 21786 20767 21788
rect 20791 21786 20847 21788
rect 20551 21734 20597 21786
rect 20597 21734 20607 21786
rect 20631 21734 20661 21786
rect 20661 21734 20673 21786
rect 20673 21734 20687 21786
rect 20711 21734 20725 21786
rect 20725 21734 20737 21786
rect 20737 21734 20767 21786
rect 20791 21734 20801 21786
rect 20801 21734 20847 21786
rect 20551 21732 20607 21734
rect 20631 21732 20687 21734
rect 20711 21732 20767 21734
rect 20791 21732 20847 21734
rect 19430 20848 19486 20904
rect 18102 19066 18158 19068
rect 18182 19066 18238 19068
rect 18262 19066 18318 19068
rect 18342 19066 18398 19068
rect 18102 19014 18148 19066
rect 18148 19014 18158 19066
rect 18182 19014 18212 19066
rect 18212 19014 18224 19066
rect 18224 19014 18238 19066
rect 18262 19014 18276 19066
rect 18276 19014 18288 19066
rect 18288 19014 18318 19066
rect 18342 19014 18352 19066
rect 18352 19014 18398 19066
rect 18102 19012 18158 19014
rect 18182 19012 18238 19014
rect 18262 19012 18318 19014
rect 18342 19012 18398 19014
rect 15652 13082 15708 13084
rect 15732 13082 15788 13084
rect 15812 13082 15868 13084
rect 15892 13082 15948 13084
rect 15652 13030 15698 13082
rect 15698 13030 15708 13082
rect 15732 13030 15762 13082
rect 15762 13030 15774 13082
rect 15774 13030 15788 13082
rect 15812 13030 15826 13082
rect 15826 13030 15838 13082
rect 15838 13030 15868 13082
rect 15892 13030 15902 13082
rect 15902 13030 15948 13082
rect 15652 13028 15708 13030
rect 15732 13028 15788 13030
rect 15812 13028 15868 13030
rect 15892 13028 15948 13030
rect 15652 11994 15708 11996
rect 15732 11994 15788 11996
rect 15812 11994 15868 11996
rect 15892 11994 15948 11996
rect 15652 11942 15698 11994
rect 15698 11942 15708 11994
rect 15732 11942 15762 11994
rect 15762 11942 15774 11994
rect 15774 11942 15788 11994
rect 15812 11942 15826 11994
rect 15826 11942 15838 11994
rect 15838 11942 15868 11994
rect 15892 11942 15902 11994
rect 15902 11942 15948 11994
rect 15652 11940 15708 11942
rect 15732 11940 15788 11942
rect 15812 11940 15868 11942
rect 15892 11940 15948 11942
rect 15652 10906 15708 10908
rect 15732 10906 15788 10908
rect 15812 10906 15868 10908
rect 15892 10906 15948 10908
rect 15652 10854 15698 10906
rect 15698 10854 15708 10906
rect 15732 10854 15762 10906
rect 15762 10854 15774 10906
rect 15774 10854 15788 10906
rect 15812 10854 15826 10906
rect 15826 10854 15838 10906
rect 15838 10854 15868 10906
rect 15892 10854 15902 10906
rect 15902 10854 15948 10906
rect 15652 10852 15708 10854
rect 15732 10852 15788 10854
rect 15812 10852 15868 10854
rect 15892 10852 15948 10854
rect 15652 9818 15708 9820
rect 15732 9818 15788 9820
rect 15812 9818 15868 9820
rect 15892 9818 15948 9820
rect 15652 9766 15698 9818
rect 15698 9766 15708 9818
rect 15732 9766 15762 9818
rect 15762 9766 15774 9818
rect 15774 9766 15788 9818
rect 15812 9766 15826 9818
rect 15826 9766 15838 9818
rect 15838 9766 15868 9818
rect 15892 9766 15902 9818
rect 15902 9766 15948 9818
rect 15652 9764 15708 9766
rect 15732 9764 15788 9766
rect 15812 9764 15868 9766
rect 15892 9764 15948 9766
rect 15652 8730 15708 8732
rect 15732 8730 15788 8732
rect 15812 8730 15868 8732
rect 15892 8730 15948 8732
rect 15652 8678 15698 8730
rect 15698 8678 15708 8730
rect 15732 8678 15762 8730
rect 15762 8678 15774 8730
rect 15774 8678 15788 8730
rect 15812 8678 15826 8730
rect 15826 8678 15838 8730
rect 15838 8678 15868 8730
rect 15892 8678 15902 8730
rect 15902 8678 15948 8730
rect 15652 8676 15708 8678
rect 15732 8676 15788 8678
rect 15812 8676 15868 8678
rect 15892 8676 15948 8678
rect 15652 7642 15708 7644
rect 15732 7642 15788 7644
rect 15812 7642 15868 7644
rect 15892 7642 15948 7644
rect 15652 7590 15698 7642
rect 15698 7590 15708 7642
rect 15732 7590 15762 7642
rect 15762 7590 15774 7642
rect 15774 7590 15788 7642
rect 15812 7590 15826 7642
rect 15826 7590 15838 7642
rect 15838 7590 15868 7642
rect 15892 7590 15902 7642
rect 15902 7590 15948 7642
rect 15652 7588 15708 7590
rect 15732 7588 15788 7590
rect 15812 7588 15868 7590
rect 15892 7588 15948 7590
rect 15652 6554 15708 6556
rect 15732 6554 15788 6556
rect 15812 6554 15868 6556
rect 15892 6554 15948 6556
rect 15652 6502 15698 6554
rect 15698 6502 15708 6554
rect 15732 6502 15762 6554
rect 15762 6502 15774 6554
rect 15774 6502 15788 6554
rect 15812 6502 15826 6554
rect 15826 6502 15838 6554
rect 15838 6502 15868 6554
rect 15892 6502 15902 6554
rect 15902 6502 15948 6554
rect 15652 6500 15708 6502
rect 15732 6500 15788 6502
rect 15812 6500 15868 6502
rect 15892 6500 15948 6502
rect 15652 5466 15708 5468
rect 15732 5466 15788 5468
rect 15812 5466 15868 5468
rect 15892 5466 15948 5468
rect 15652 5414 15698 5466
rect 15698 5414 15708 5466
rect 15732 5414 15762 5466
rect 15762 5414 15774 5466
rect 15774 5414 15788 5466
rect 15812 5414 15826 5466
rect 15826 5414 15838 5466
rect 15838 5414 15868 5466
rect 15892 5414 15902 5466
rect 15902 5414 15948 5466
rect 15652 5412 15708 5414
rect 15732 5412 15788 5414
rect 15812 5412 15868 5414
rect 15892 5412 15948 5414
rect 15652 4378 15708 4380
rect 15732 4378 15788 4380
rect 15812 4378 15868 4380
rect 15892 4378 15948 4380
rect 15652 4326 15698 4378
rect 15698 4326 15708 4378
rect 15732 4326 15762 4378
rect 15762 4326 15774 4378
rect 15774 4326 15788 4378
rect 15812 4326 15826 4378
rect 15826 4326 15838 4378
rect 15838 4326 15868 4378
rect 15892 4326 15902 4378
rect 15902 4326 15948 4378
rect 15652 4324 15708 4326
rect 15732 4324 15788 4326
rect 15812 4324 15868 4326
rect 15892 4324 15948 4326
rect 15652 3290 15708 3292
rect 15732 3290 15788 3292
rect 15812 3290 15868 3292
rect 15892 3290 15948 3292
rect 15652 3238 15698 3290
rect 15698 3238 15708 3290
rect 15732 3238 15762 3290
rect 15762 3238 15774 3290
rect 15774 3238 15788 3290
rect 15812 3238 15826 3290
rect 15826 3238 15838 3290
rect 15838 3238 15868 3290
rect 15892 3238 15902 3290
rect 15902 3238 15948 3290
rect 15652 3236 15708 3238
rect 15732 3236 15788 3238
rect 15812 3236 15868 3238
rect 15892 3236 15948 3238
rect 18102 17978 18158 17980
rect 18182 17978 18238 17980
rect 18262 17978 18318 17980
rect 18342 17978 18398 17980
rect 18102 17926 18148 17978
rect 18148 17926 18158 17978
rect 18182 17926 18212 17978
rect 18212 17926 18224 17978
rect 18224 17926 18238 17978
rect 18262 17926 18276 17978
rect 18276 17926 18288 17978
rect 18288 17926 18318 17978
rect 18342 17926 18352 17978
rect 18352 17926 18398 17978
rect 18102 17924 18158 17926
rect 18182 17924 18238 17926
rect 18262 17924 18318 17926
rect 18342 17924 18398 17926
rect 18102 16890 18158 16892
rect 18182 16890 18238 16892
rect 18262 16890 18318 16892
rect 18342 16890 18398 16892
rect 18102 16838 18148 16890
rect 18148 16838 18158 16890
rect 18182 16838 18212 16890
rect 18212 16838 18224 16890
rect 18224 16838 18238 16890
rect 18262 16838 18276 16890
rect 18276 16838 18288 16890
rect 18288 16838 18318 16890
rect 18342 16838 18352 16890
rect 18352 16838 18398 16890
rect 18102 16836 18158 16838
rect 18182 16836 18238 16838
rect 18262 16836 18318 16838
rect 18342 16836 18398 16838
rect 18102 15802 18158 15804
rect 18182 15802 18238 15804
rect 18262 15802 18318 15804
rect 18342 15802 18398 15804
rect 18102 15750 18148 15802
rect 18148 15750 18158 15802
rect 18182 15750 18212 15802
rect 18212 15750 18224 15802
rect 18224 15750 18238 15802
rect 18262 15750 18276 15802
rect 18276 15750 18288 15802
rect 18288 15750 18318 15802
rect 18342 15750 18352 15802
rect 18352 15750 18398 15802
rect 18102 15748 18158 15750
rect 18182 15748 18238 15750
rect 18262 15748 18318 15750
rect 18342 15748 18398 15750
rect 18102 14714 18158 14716
rect 18182 14714 18238 14716
rect 18262 14714 18318 14716
rect 18342 14714 18398 14716
rect 18102 14662 18148 14714
rect 18148 14662 18158 14714
rect 18182 14662 18212 14714
rect 18212 14662 18224 14714
rect 18224 14662 18238 14714
rect 18262 14662 18276 14714
rect 18276 14662 18288 14714
rect 18288 14662 18318 14714
rect 18342 14662 18352 14714
rect 18352 14662 18398 14714
rect 18102 14660 18158 14662
rect 18182 14660 18238 14662
rect 18262 14660 18318 14662
rect 18342 14660 18398 14662
rect 18102 13626 18158 13628
rect 18182 13626 18238 13628
rect 18262 13626 18318 13628
rect 18342 13626 18398 13628
rect 18102 13574 18148 13626
rect 18148 13574 18158 13626
rect 18182 13574 18212 13626
rect 18212 13574 18224 13626
rect 18224 13574 18238 13626
rect 18262 13574 18276 13626
rect 18276 13574 18288 13626
rect 18288 13574 18318 13626
rect 18342 13574 18352 13626
rect 18352 13574 18398 13626
rect 18102 13572 18158 13574
rect 18182 13572 18238 13574
rect 18262 13572 18318 13574
rect 18342 13572 18398 13574
rect 18102 12538 18158 12540
rect 18182 12538 18238 12540
rect 18262 12538 18318 12540
rect 18342 12538 18398 12540
rect 18102 12486 18148 12538
rect 18148 12486 18158 12538
rect 18182 12486 18212 12538
rect 18212 12486 18224 12538
rect 18224 12486 18238 12538
rect 18262 12486 18276 12538
rect 18276 12486 18288 12538
rect 18288 12486 18318 12538
rect 18342 12486 18352 12538
rect 18352 12486 18398 12538
rect 18102 12484 18158 12486
rect 18182 12484 18238 12486
rect 18262 12484 18318 12486
rect 18342 12484 18398 12486
rect 18102 11450 18158 11452
rect 18182 11450 18238 11452
rect 18262 11450 18318 11452
rect 18342 11450 18398 11452
rect 18102 11398 18148 11450
rect 18148 11398 18158 11450
rect 18182 11398 18212 11450
rect 18212 11398 18224 11450
rect 18224 11398 18238 11450
rect 18262 11398 18276 11450
rect 18276 11398 18288 11450
rect 18288 11398 18318 11450
rect 18342 11398 18352 11450
rect 18352 11398 18398 11450
rect 18102 11396 18158 11398
rect 18182 11396 18238 11398
rect 18262 11396 18318 11398
rect 18342 11396 18398 11398
rect 18102 10362 18158 10364
rect 18182 10362 18238 10364
rect 18262 10362 18318 10364
rect 18342 10362 18398 10364
rect 18102 10310 18148 10362
rect 18148 10310 18158 10362
rect 18182 10310 18212 10362
rect 18212 10310 18224 10362
rect 18224 10310 18238 10362
rect 18262 10310 18276 10362
rect 18276 10310 18288 10362
rect 18288 10310 18318 10362
rect 18342 10310 18352 10362
rect 18352 10310 18398 10362
rect 18102 10308 18158 10310
rect 18182 10308 18238 10310
rect 18262 10308 18318 10310
rect 18342 10308 18398 10310
rect 18102 9274 18158 9276
rect 18182 9274 18238 9276
rect 18262 9274 18318 9276
rect 18342 9274 18398 9276
rect 18102 9222 18148 9274
rect 18148 9222 18158 9274
rect 18182 9222 18212 9274
rect 18212 9222 18224 9274
rect 18224 9222 18238 9274
rect 18262 9222 18276 9274
rect 18276 9222 18288 9274
rect 18288 9222 18318 9274
rect 18342 9222 18352 9274
rect 18352 9222 18398 9274
rect 18102 9220 18158 9222
rect 18182 9220 18238 9222
rect 18262 9220 18318 9222
rect 18342 9220 18398 9222
rect 18102 8186 18158 8188
rect 18182 8186 18238 8188
rect 18262 8186 18318 8188
rect 18342 8186 18398 8188
rect 18102 8134 18148 8186
rect 18148 8134 18158 8186
rect 18182 8134 18212 8186
rect 18212 8134 18224 8186
rect 18224 8134 18238 8186
rect 18262 8134 18276 8186
rect 18276 8134 18288 8186
rect 18288 8134 18318 8186
rect 18342 8134 18352 8186
rect 18352 8134 18398 8186
rect 18102 8132 18158 8134
rect 18182 8132 18238 8134
rect 18262 8132 18318 8134
rect 18342 8132 18398 8134
rect 18102 7098 18158 7100
rect 18182 7098 18238 7100
rect 18262 7098 18318 7100
rect 18342 7098 18398 7100
rect 18102 7046 18148 7098
rect 18148 7046 18158 7098
rect 18182 7046 18212 7098
rect 18212 7046 18224 7098
rect 18224 7046 18238 7098
rect 18262 7046 18276 7098
rect 18276 7046 18288 7098
rect 18288 7046 18318 7098
rect 18342 7046 18352 7098
rect 18352 7046 18398 7098
rect 18102 7044 18158 7046
rect 18182 7044 18238 7046
rect 18262 7044 18318 7046
rect 18342 7044 18398 7046
rect 18102 6010 18158 6012
rect 18182 6010 18238 6012
rect 18262 6010 18318 6012
rect 18342 6010 18398 6012
rect 18102 5958 18148 6010
rect 18148 5958 18158 6010
rect 18182 5958 18212 6010
rect 18212 5958 18224 6010
rect 18224 5958 18238 6010
rect 18262 5958 18276 6010
rect 18276 5958 18288 6010
rect 18288 5958 18318 6010
rect 18342 5958 18352 6010
rect 18352 5958 18398 6010
rect 18102 5956 18158 5958
rect 18182 5956 18238 5958
rect 18262 5956 18318 5958
rect 18342 5956 18398 5958
rect 18102 4922 18158 4924
rect 18182 4922 18238 4924
rect 18262 4922 18318 4924
rect 18342 4922 18398 4924
rect 18102 4870 18148 4922
rect 18148 4870 18158 4922
rect 18182 4870 18212 4922
rect 18212 4870 18224 4922
rect 18224 4870 18238 4922
rect 18262 4870 18276 4922
rect 18276 4870 18288 4922
rect 18288 4870 18318 4922
rect 18342 4870 18352 4922
rect 18352 4870 18398 4922
rect 18102 4868 18158 4870
rect 18182 4868 18238 4870
rect 18262 4868 18318 4870
rect 18342 4868 18398 4870
rect 18102 3834 18158 3836
rect 18182 3834 18238 3836
rect 18262 3834 18318 3836
rect 18342 3834 18398 3836
rect 18102 3782 18148 3834
rect 18148 3782 18158 3834
rect 18182 3782 18212 3834
rect 18212 3782 18224 3834
rect 18224 3782 18238 3834
rect 18262 3782 18276 3834
rect 18276 3782 18288 3834
rect 18288 3782 18318 3834
rect 18342 3782 18352 3834
rect 18352 3782 18398 3834
rect 18102 3780 18158 3782
rect 18182 3780 18238 3782
rect 18262 3780 18318 3782
rect 18342 3780 18398 3782
rect 18102 2746 18158 2748
rect 18182 2746 18238 2748
rect 18262 2746 18318 2748
rect 18342 2746 18398 2748
rect 18102 2694 18148 2746
rect 18148 2694 18158 2746
rect 18182 2694 18212 2746
rect 18212 2694 18224 2746
rect 18224 2694 18238 2746
rect 18262 2694 18276 2746
rect 18276 2694 18288 2746
rect 18288 2694 18318 2746
rect 18342 2694 18352 2746
rect 18352 2694 18398 2746
rect 18102 2692 18158 2694
rect 18182 2692 18238 2694
rect 18262 2692 18318 2694
rect 18342 2692 18398 2694
rect 5854 2202 5910 2204
rect 5934 2202 5990 2204
rect 6014 2202 6070 2204
rect 6094 2202 6150 2204
rect 5854 2150 5900 2202
rect 5900 2150 5910 2202
rect 5934 2150 5964 2202
rect 5964 2150 5976 2202
rect 5976 2150 5990 2202
rect 6014 2150 6028 2202
rect 6028 2150 6040 2202
rect 6040 2150 6070 2202
rect 6094 2150 6104 2202
rect 6104 2150 6150 2202
rect 5854 2148 5910 2150
rect 5934 2148 5990 2150
rect 6014 2148 6070 2150
rect 6094 2148 6150 2150
rect 10753 2202 10809 2204
rect 10833 2202 10889 2204
rect 10913 2202 10969 2204
rect 10993 2202 11049 2204
rect 10753 2150 10799 2202
rect 10799 2150 10809 2202
rect 10833 2150 10863 2202
rect 10863 2150 10875 2202
rect 10875 2150 10889 2202
rect 10913 2150 10927 2202
rect 10927 2150 10939 2202
rect 10939 2150 10969 2202
rect 10993 2150 11003 2202
rect 11003 2150 11049 2202
rect 10753 2148 10809 2150
rect 10833 2148 10889 2150
rect 10913 2148 10969 2150
rect 10993 2148 11049 2150
rect 15652 2202 15708 2204
rect 15732 2202 15788 2204
rect 15812 2202 15868 2204
rect 15892 2202 15948 2204
rect 15652 2150 15698 2202
rect 15698 2150 15708 2202
rect 15732 2150 15762 2202
rect 15762 2150 15774 2202
rect 15774 2150 15788 2202
rect 15812 2150 15826 2202
rect 15826 2150 15838 2202
rect 15838 2150 15868 2202
rect 15892 2150 15902 2202
rect 15902 2150 15948 2202
rect 15652 2148 15708 2150
rect 15732 2148 15788 2150
rect 15812 2148 15868 2150
rect 15892 2148 15948 2150
rect 20551 20698 20607 20700
rect 20631 20698 20687 20700
rect 20711 20698 20767 20700
rect 20791 20698 20847 20700
rect 20551 20646 20597 20698
rect 20597 20646 20607 20698
rect 20631 20646 20661 20698
rect 20661 20646 20673 20698
rect 20673 20646 20687 20698
rect 20711 20646 20725 20698
rect 20725 20646 20737 20698
rect 20737 20646 20767 20698
rect 20791 20646 20801 20698
rect 20801 20646 20847 20698
rect 20551 20644 20607 20646
rect 20631 20644 20687 20646
rect 20711 20644 20767 20646
rect 20791 20644 20847 20646
rect 20551 19610 20607 19612
rect 20631 19610 20687 19612
rect 20711 19610 20767 19612
rect 20791 19610 20847 19612
rect 20551 19558 20597 19610
rect 20597 19558 20607 19610
rect 20631 19558 20661 19610
rect 20661 19558 20673 19610
rect 20673 19558 20687 19610
rect 20711 19558 20725 19610
rect 20725 19558 20737 19610
rect 20737 19558 20767 19610
rect 20791 19558 20801 19610
rect 20801 19558 20847 19610
rect 20551 19556 20607 19558
rect 20631 19556 20687 19558
rect 20711 19556 20767 19558
rect 20791 19556 20847 19558
rect 20074 19080 20130 19136
rect 19982 17856 20038 17912
rect 19982 15544 20038 15600
rect 20551 18522 20607 18524
rect 20631 18522 20687 18524
rect 20711 18522 20767 18524
rect 20791 18522 20847 18524
rect 20551 18470 20597 18522
rect 20597 18470 20607 18522
rect 20631 18470 20661 18522
rect 20661 18470 20673 18522
rect 20673 18470 20687 18522
rect 20711 18470 20725 18522
rect 20725 18470 20737 18522
rect 20737 18470 20767 18522
rect 20791 18470 20801 18522
rect 20801 18470 20847 18522
rect 20551 18468 20607 18470
rect 20631 18468 20687 18470
rect 20711 18468 20767 18470
rect 20791 18468 20847 18470
rect 20551 17434 20607 17436
rect 20631 17434 20687 17436
rect 20711 17434 20767 17436
rect 20791 17434 20847 17436
rect 20551 17382 20597 17434
rect 20597 17382 20607 17434
rect 20631 17382 20661 17434
rect 20661 17382 20673 17434
rect 20673 17382 20687 17434
rect 20711 17382 20725 17434
rect 20725 17382 20737 17434
rect 20737 17382 20767 17434
rect 20791 17382 20801 17434
rect 20801 17382 20847 17434
rect 20551 17380 20607 17382
rect 20631 17380 20687 17382
rect 20711 17380 20767 17382
rect 20791 17380 20847 17382
rect 20551 16346 20607 16348
rect 20631 16346 20687 16348
rect 20711 16346 20767 16348
rect 20791 16346 20847 16348
rect 20551 16294 20597 16346
rect 20597 16294 20607 16346
rect 20631 16294 20661 16346
rect 20661 16294 20673 16346
rect 20673 16294 20687 16346
rect 20711 16294 20725 16346
rect 20725 16294 20737 16346
rect 20737 16294 20767 16346
rect 20791 16294 20801 16346
rect 20801 16294 20847 16346
rect 20551 16292 20607 16294
rect 20631 16292 20687 16294
rect 20711 16292 20767 16294
rect 20791 16292 20847 16294
rect 20551 15258 20607 15260
rect 20631 15258 20687 15260
rect 20711 15258 20767 15260
rect 20791 15258 20847 15260
rect 20551 15206 20597 15258
rect 20597 15206 20607 15258
rect 20631 15206 20661 15258
rect 20661 15206 20673 15258
rect 20673 15206 20687 15258
rect 20711 15206 20725 15258
rect 20725 15206 20737 15258
rect 20737 15206 20767 15258
rect 20791 15206 20801 15258
rect 20801 15206 20847 15258
rect 20551 15204 20607 15206
rect 20631 15204 20687 15206
rect 20711 15204 20767 15206
rect 20791 15204 20847 15206
rect 20551 14170 20607 14172
rect 20631 14170 20687 14172
rect 20711 14170 20767 14172
rect 20791 14170 20847 14172
rect 20551 14118 20597 14170
rect 20597 14118 20607 14170
rect 20631 14118 20661 14170
rect 20661 14118 20673 14170
rect 20673 14118 20687 14170
rect 20711 14118 20725 14170
rect 20725 14118 20737 14170
rect 20737 14118 20767 14170
rect 20791 14118 20801 14170
rect 20801 14118 20847 14170
rect 20551 14116 20607 14118
rect 20631 14116 20687 14118
rect 20711 14116 20767 14118
rect 20791 14116 20847 14118
rect 19982 13776 20038 13832
rect 20551 13082 20607 13084
rect 20631 13082 20687 13084
rect 20711 13082 20767 13084
rect 20791 13082 20847 13084
rect 20551 13030 20597 13082
rect 20597 13030 20607 13082
rect 20631 13030 20661 13082
rect 20661 13030 20673 13082
rect 20673 13030 20687 13082
rect 20711 13030 20725 13082
rect 20725 13030 20737 13082
rect 20737 13030 20767 13082
rect 20791 13030 20801 13082
rect 20801 13030 20847 13082
rect 20551 13028 20607 13030
rect 20631 13028 20687 13030
rect 20711 13028 20767 13030
rect 20791 13028 20847 13030
rect 19982 12316 19984 12336
rect 19984 12316 20036 12336
rect 20036 12316 20038 12336
rect 19982 12280 20038 12316
rect 20551 11994 20607 11996
rect 20631 11994 20687 11996
rect 20711 11994 20767 11996
rect 20791 11994 20847 11996
rect 20551 11942 20597 11994
rect 20597 11942 20607 11994
rect 20631 11942 20661 11994
rect 20661 11942 20673 11994
rect 20673 11942 20687 11994
rect 20711 11942 20725 11994
rect 20725 11942 20737 11994
rect 20737 11942 20767 11994
rect 20791 11942 20801 11994
rect 20801 11942 20847 11994
rect 20551 11940 20607 11942
rect 20631 11940 20687 11942
rect 20711 11940 20767 11942
rect 20791 11940 20847 11942
rect 20551 10906 20607 10908
rect 20631 10906 20687 10908
rect 20711 10906 20767 10908
rect 20791 10906 20847 10908
rect 20551 10854 20597 10906
rect 20597 10854 20607 10906
rect 20631 10854 20661 10906
rect 20661 10854 20673 10906
rect 20673 10854 20687 10906
rect 20711 10854 20725 10906
rect 20725 10854 20737 10906
rect 20737 10854 20767 10906
rect 20791 10854 20801 10906
rect 20801 10854 20847 10906
rect 20551 10852 20607 10854
rect 20631 10852 20687 10854
rect 20711 10852 20767 10854
rect 20791 10852 20847 10854
rect 19982 10260 20038 10296
rect 19982 10240 19984 10260
rect 19984 10240 20036 10260
rect 20036 10240 20038 10260
rect 20551 9818 20607 9820
rect 20631 9818 20687 9820
rect 20711 9818 20767 9820
rect 20791 9818 20847 9820
rect 20551 9766 20597 9818
rect 20597 9766 20607 9818
rect 20631 9766 20661 9818
rect 20661 9766 20673 9818
rect 20673 9766 20687 9818
rect 20711 9766 20725 9818
rect 20725 9766 20737 9818
rect 20737 9766 20767 9818
rect 20791 9766 20801 9818
rect 20801 9766 20847 9818
rect 20551 9764 20607 9766
rect 20631 9764 20687 9766
rect 20711 9764 20767 9766
rect 20791 9764 20847 9766
rect 19982 8472 20038 8528
rect 20551 8730 20607 8732
rect 20631 8730 20687 8732
rect 20711 8730 20767 8732
rect 20791 8730 20847 8732
rect 20551 8678 20597 8730
rect 20597 8678 20607 8730
rect 20631 8678 20661 8730
rect 20661 8678 20673 8730
rect 20673 8678 20687 8730
rect 20711 8678 20725 8730
rect 20725 8678 20737 8730
rect 20737 8678 20767 8730
rect 20791 8678 20801 8730
rect 20801 8678 20847 8730
rect 20551 8676 20607 8678
rect 20631 8676 20687 8678
rect 20711 8676 20767 8678
rect 20791 8676 20847 8678
rect 20551 7642 20607 7644
rect 20631 7642 20687 7644
rect 20711 7642 20767 7644
rect 20791 7642 20847 7644
rect 20551 7590 20597 7642
rect 20597 7590 20607 7642
rect 20631 7590 20661 7642
rect 20661 7590 20673 7642
rect 20673 7590 20687 7642
rect 20711 7590 20725 7642
rect 20725 7590 20737 7642
rect 20737 7590 20767 7642
rect 20791 7590 20801 7642
rect 20801 7590 20847 7642
rect 20551 7588 20607 7590
rect 20631 7588 20687 7590
rect 20711 7588 20767 7590
rect 20791 7588 20847 7590
rect 19982 6704 20038 6760
rect 20551 6554 20607 6556
rect 20631 6554 20687 6556
rect 20711 6554 20767 6556
rect 20791 6554 20847 6556
rect 20551 6502 20597 6554
rect 20597 6502 20607 6554
rect 20631 6502 20661 6554
rect 20661 6502 20673 6554
rect 20673 6502 20687 6554
rect 20711 6502 20725 6554
rect 20725 6502 20737 6554
rect 20737 6502 20767 6554
rect 20791 6502 20801 6554
rect 20801 6502 20847 6554
rect 20551 6500 20607 6502
rect 20631 6500 20687 6502
rect 20711 6500 20767 6502
rect 20791 6500 20847 6502
rect 20551 5466 20607 5468
rect 20631 5466 20687 5468
rect 20711 5466 20767 5468
rect 20791 5466 20847 5468
rect 20551 5414 20597 5466
rect 20597 5414 20607 5466
rect 20631 5414 20661 5466
rect 20661 5414 20673 5466
rect 20673 5414 20687 5466
rect 20711 5414 20725 5466
rect 20725 5414 20737 5466
rect 20737 5414 20767 5466
rect 20791 5414 20801 5466
rect 20801 5414 20847 5466
rect 20551 5412 20607 5414
rect 20631 5412 20687 5414
rect 20711 5412 20767 5414
rect 20791 5412 20847 5414
rect 20074 4972 20076 4992
rect 20076 4972 20128 4992
rect 20128 4972 20130 4992
rect 20074 4936 20130 4972
rect 20551 4378 20607 4380
rect 20631 4378 20687 4380
rect 20711 4378 20767 4380
rect 20791 4378 20847 4380
rect 20551 4326 20597 4378
rect 20597 4326 20607 4378
rect 20631 4326 20661 4378
rect 20661 4326 20673 4378
rect 20673 4326 20687 4378
rect 20711 4326 20725 4378
rect 20725 4326 20737 4378
rect 20737 4326 20767 4378
rect 20791 4326 20801 4378
rect 20801 4326 20847 4378
rect 20551 4324 20607 4326
rect 20631 4324 20687 4326
rect 20711 4324 20767 4326
rect 20791 4324 20847 4326
rect 20074 3440 20130 3496
rect 20551 3290 20607 3292
rect 20631 3290 20687 3292
rect 20711 3290 20767 3292
rect 20791 3290 20847 3292
rect 20551 3238 20597 3290
rect 20597 3238 20607 3290
rect 20631 3238 20661 3290
rect 20661 3238 20673 3290
rect 20673 3238 20687 3290
rect 20711 3238 20725 3290
rect 20725 3238 20737 3290
rect 20737 3238 20767 3290
rect 20791 3238 20801 3290
rect 20801 3238 20847 3290
rect 20551 3236 20607 3238
rect 20631 3236 20687 3238
rect 20711 3236 20767 3238
rect 20791 3236 20847 3238
rect 19154 1400 19210 1456
rect 20551 2202 20607 2204
rect 20631 2202 20687 2204
rect 20711 2202 20767 2204
rect 20791 2202 20847 2204
rect 20551 2150 20597 2202
rect 20597 2150 20607 2202
rect 20631 2150 20661 2202
rect 20661 2150 20673 2202
rect 20673 2150 20687 2202
rect 20711 2150 20725 2202
rect 20725 2150 20737 2202
rect 20737 2150 20767 2202
rect 20791 2150 20801 2202
rect 20801 2150 20847 2202
rect 20551 2148 20607 2150
rect 20631 2148 20687 2150
rect 20711 2148 20767 2150
rect 20791 2148 20847 2150
<< metal3 >>
rect 16481 22674 16547 22677
rect 21061 22674 21861 22704
rect 16481 22672 21861 22674
rect 16481 22616 16486 22672
rect 16542 22616 21861 22672
rect 16481 22614 21861 22616
rect 16481 22611 16547 22614
rect 21061 22584 21861 22614
rect 0 21858 800 21888
rect 1669 21858 1735 21861
rect 0 21856 1735 21858
rect 0 21800 1674 21856
rect 1730 21800 1735 21856
rect 0 21798 1735 21800
rect 0 21768 800 21798
rect 1669 21795 1735 21798
rect 5844 21792 6160 21793
rect 5844 21728 5850 21792
rect 5914 21728 5930 21792
rect 5994 21728 6010 21792
rect 6074 21728 6090 21792
rect 6154 21728 6160 21792
rect 5844 21727 6160 21728
rect 10743 21792 11059 21793
rect 10743 21728 10749 21792
rect 10813 21728 10829 21792
rect 10893 21728 10909 21792
rect 10973 21728 10989 21792
rect 11053 21728 11059 21792
rect 10743 21727 11059 21728
rect 15642 21792 15958 21793
rect 15642 21728 15648 21792
rect 15712 21728 15728 21792
rect 15792 21728 15808 21792
rect 15872 21728 15888 21792
rect 15952 21728 15958 21792
rect 15642 21727 15958 21728
rect 20541 21792 20857 21793
rect 20541 21728 20547 21792
rect 20611 21728 20627 21792
rect 20691 21728 20707 21792
rect 20771 21728 20787 21792
rect 20851 21728 20857 21792
rect 20541 21727 20857 21728
rect 3395 21248 3711 21249
rect 3395 21184 3401 21248
rect 3465 21184 3481 21248
rect 3545 21184 3561 21248
rect 3625 21184 3641 21248
rect 3705 21184 3711 21248
rect 3395 21183 3711 21184
rect 8294 21248 8610 21249
rect 8294 21184 8300 21248
rect 8364 21184 8380 21248
rect 8444 21184 8460 21248
rect 8524 21184 8540 21248
rect 8604 21184 8610 21248
rect 8294 21183 8610 21184
rect 13193 21248 13509 21249
rect 13193 21184 13199 21248
rect 13263 21184 13279 21248
rect 13343 21184 13359 21248
rect 13423 21184 13439 21248
rect 13503 21184 13509 21248
rect 13193 21183 13509 21184
rect 18092 21248 18408 21249
rect 18092 21184 18098 21248
rect 18162 21184 18178 21248
rect 18242 21184 18258 21248
rect 18322 21184 18338 21248
rect 18402 21184 18408 21248
rect 18092 21183 18408 21184
rect 19425 20906 19491 20909
rect 21061 20906 21861 20936
rect 19425 20904 21861 20906
rect 19425 20848 19430 20904
rect 19486 20848 21861 20904
rect 19425 20846 21861 20848
rect 19425 20843 19491 20846
rect 21061 20816 21861 20846
rect 5844 20704 6160 20705
rect 5844 20640 5850 20704
rect 5914 20640 5930 20704
rect 5994 20640 6010 20704
rect 6074 20640 6090 20704
rect 6154 20640 6160 20704
rect 5844 20639 6160 20640
rect 10743 20704 11059 20705
rect 10743 20640 10749 20704
rect 10813 20640 10829 20704
rect 10893 20640 10909 20704
rect 10973 20640 10989 20704
rect 11053 20640 11059 20704
rect 10743 20639 11059 20640
rect 15642 20704 15958 20705
rect 15642 20640 15648 20704
rect 15712 20640 15728 20704
rect 15792 20640 15808 20704
rect 15872 20640 15888 20704
rect 15952 20640 15958 20704
rect 15642 20639 15958 20640
rect 20541 20704 20857 20705
rect 20541 20640 20547 20704
rect 20611 20640 20627 20704
rect 20691 20640 20707 20704
rect 20771 20640 20787 20704
rect 20851 20640 20857 20704
rect 20541 20639 20857 20640
rect 3395 20160 3711 20161
rect 3395 20096 3401 20160
rect 3465 20096 3481 20160
rect 3545 20096 3561 20160
rect 3625 20096 3641 20160
rect 3705 20096 3711 20160
rect 3395 20095 3711 20096
rect 8294 20160 8610 20161
rect 8294 20096 8300 20160
rect 8364 20096 8380 20160
rect 8444 20096 8460 20160
rect 8524 20096 8540 20160
rect 8604 20096 8610 20160
rect 8294 20095 8610 20096
rect 13193 20160 13509 20161
rect 13193 20096 13199 20160
rect 13263 20096 13279 20160
rect 13343 20096 13359 20160
rect 13423 20096 13439 20160
rect 13503 20096 13509 20160
rect 13193 20095 13509 20096
rect 18092 20160 18408 20161
rect 18092 20096 18098 20160
rect 18162 20096 18178 20160
rect 18242 20096 18258 20160
rect 18322 20096 18338 20160
rect 18402 20096 18408 20160
rect 18092 20095 18408 20096
rect 5844 19616 6160 19617
rect 5844 19552 5850 19616
rect 5914 19552 5930 19616
rect 5994 19552 6010 19616
rect 6074 19552 6090 19616
rect 6154 19552 6160 19616
rect 5844 19551 6160 19552
rect 10743 19616 11059 19617
rect 10743 19552 10749 19616
rect 10813 19552 10829 19616
rect 10893 19552 10909 19616
rect 10973 19552 10989 19616
rect 11053 19552 11059 19616
rect 10743 19551 11059 19552
rect 15642 19616 15958 19617
rect 15642 19552 15648 19616
rect 15712 19552 15728 19616
rect 15792 19552 15808 19616
rect 15872 19552 15888 19616
rect 15952 19552 15958 19616
rect 15642 19551 15958 19552
rect 20541 19616 20857 19617
rect 20541 19552 20547 19616
rect 20611 19552 20627 19616
rect 20691 19552 20707 19616
rect 20771 19552 20787 19616
rect 20851 19552 20857 19616
rect 20541 19551 20857 19552
rect 20069 19138 20135 19141
rect 21061 19138 21861 19168
rect 20069 19136 21861 19138
rect 20069 19080 20074 19136
rect 20130 19080 21861 19136
rect 20069 19078 21861 19080
rect 20069 19075 20135 19078
rect 3395 19072 3711 19073
rect 3395 19008 3401 19072
rect 3465 19008 3481 19072
rect 3545 19008 3561 19072
rect 3625 19008 3641 19072
rect 3705 19008 3711 19072
rect 3395 19007 3711 19008
rect 8294 19072 8610 19073
rect 8294 19008 8300 19072
rect 8364 19008 8380 19072
rect 8444 19008 8460 19072
rect 8524 19008 8540 19072
rect 8604 19008 8610 19072
rect 8294 19007 8610 19008
rect 13193 19072 13509 19073
rect 13193 19008 13199 19072
rect 13263 19008 13279 19072
rect 13343 19008 13359 19072
rect 13423 19008 13439 19072
rect 13503 19008 13509 19072
rect 13193 19007 13509 19008
rect 18092 19072 18408 19073
rect 18092 19008 18098 19072
rect 18162 19008 18178 19072
rect 18242 19008 18258 19072
rect 18322 19008 18338 19072
rect 18402 19008 18408 19072
rect 21061 19048 21861 19078
rect 18092 19007 18408 19008
rect 800 18540 1480 18560
rect 800 18460 1120 18540
rect 1470 18460 1480 18540
rect 5844 18528 6160 18529
rect 5844 18464 5850 18528
rect 5914 18464 5930 18528
rect 5994 18464 6010 18528
rect 6074 18464 6090 18528
rect 6154 18464 6160 18528
rect 5844 18463 6160 18464
rect 10743 18528 11059 18529
rect 10743 18464 10749 18528
rect 10813 18464 10829 18528
rect 10893 18464 10909 18528
rect 10973 18464 10989 18528
rect 11053 18464 11059 18528
rect 10743 18463 11059 18464
rect 15642 18528 15958 18529
rect 15642 18464 15648 18528
rect 15712 18464 15728 18528
rect 15792 18464 15808 18528
rect 15872 18464 15888 18528
rect 15952 18464 15958 18528
rect 15642 18463 15958 18464
rect 20541 18528 20857 18529
rect 20541 18464 20547 18528
rect 20611 18464 20627 18528
rect 20691 18464 20707 18528
rect 20771 18464 20787 18528
rect 20851 18464 20857 18528
rect 20541 18463 20857 18464
rect 800 18440 1480 18460
rect 800 17944 920 18440
rect 0 17840 920 17944
rect 3395 17984 3711 17985
rect 3395 17920 3401 17984
rect 3465 17920 3481 17984
rect 3545 17920 3561 17984
rect 3625 17920 3641 17984
rect 3705 17920 3711 17984
rect 3395 17919 3711 17920
rect 8294 17984 8610 17985
rect 8294 17920 8300 17984
rect 8364 17920 8380 17984
rect 8444 17920 8460 17984
rect 8524 17920 8540 17984
rect 8604 17920 8610 17984
rect 8294 17919 8610 17920
rect 13193 17984 13509 17985
rect 13193 17920 13199 17984
rect 13263 17920 13279 17984
rect 13343 17920 13359 17984
rect 13423 17920 13439 17984
rect 13503 17920 13509 17984
rect 13193 17919 13509 17920
rect 18092 17984 18408 17985
rect 18092 17920 18098 17984
rect 18162 17920 18178 17984
rect 18242 17920 18258 17984
rect 18322 17920 18338 17984
rect 18402 17920 18408 17984
rect 18092 17919 18408 17920
rect 19977 17914 20043 17917
rect 19977 17912 21282 17914
rect 19977 17856 19982 17912
rect 20038 17856 21282 17912
rect 19977 17854 21282 17856
rect 19977 17851 20043 17854
rect 0 17824 800 17840
rect 5844 17440 6160 17441
rect 5844 17376 5850 17440
rect 5914 17376 5930 17440
rect 5994 17376 6010 17440
rect 6074 17376 6090 17440
rect 6154 17376 6160 17440
rect 5844 17375 6160 17376
rect 10743 17440 11059 17441
rect 10743 17376 10749 17440
rect 10813 17376 10829 17440
rect 10893 17376 10909 17440
rect 10973 17376 10989 17440
rect 11053 17376 11059 17440
rect 10743 17375 11059 17376
rect 15642 17440 15958 17441
rect 15642 17376 15648 17440
rect 15712 17376 15728 17440
rect 15792 17376 15808 17440
rect 15872 17376 15888 17440
rect 15952 17376 15958 17440
rect 15642 17375 15958 17376
rect 20541 17440 20857 17441
rect 20541 17376 20547 17440
rect 20611 17376 20627 17440
rect 20691 17376 20707 17440
rect 20771 17376 20787 17440
rect 20851 17376 20857 17440
rect 21222 17400 21282 17854
rect 20541 17375 20857 17376
rect 21061 17280 21861 17400
rect 3395 16896 3711 16897
rect 3395 16832 3401 16896
rect 3465 16832 3481 16896
rect 3545 16832 3561 16896
rect 3625 16832 3641 16896
rect 3705 16832 3711 16896
rect 3395 16831 3711 16832
rect 8294 16896 8610 16897
rect 8294 16832 8300 16896
rect 8364 16832 8380 16896
rect 8444 16832 8460 16896
rect 8524 16832 8540 16896
rect 8604 16832 8610 16896
rect 8294 16831 8610 16832
rect 13193 16896 13509 16897
rect 13193 16832 13199 16896
rect 13263 16832 13279 16896
rect 13343 16832 13359 16896
rect 13423 16832 13439 16896
rect 13503 16832 13509 16896
rect 13193 16831 13509 16832
rect 18092 16896 18408 16897
rect 18092 16832 18098 16896
rect 18162 16832 18178 16896
rect 18242 16832 18258 16896
rect 18322 16832 18338 16896
rect 18402 16832 18408 16896
rect 18092 16831 18408 16832
rect 5844 16352 6160 16353
rect 5844 16288 5850 16352
rect 5914 16288 5930 16352
rect 5994 16288 6010 16352
rect 6074 16288 6090 16352
rect 6154 16288 6160 16352
rect 5844 16287 6160 16288
rect 10743 16352 11059 16353
rect 10743 16288 10749 16352
rect 10813 16288 10829 16352
rect 10893 16288 10909 16352
rect 10973 16288 10989 16352
rect 11053 16288 11059 16352
rect 10743 16287 11059 16288
rect 15642 16352 15958 16353
rect 15642 16288 15648 16352
rect 15712 16288 15728 16352
rect 15792 16288 15808 16352
rect 15872 16288 15888 16352
rect 15952 16288 15958 16352
rect 15642 16287 15958 16288
rect 20541 16352 20857 16353
rect 20541 16288 20547 16352
rect 20611 16288 20627 16352
rect 20691 16288 20707 16352
rect 20771 16288 20787 16352
rect 20851 16288 20857 16352
rect 20541 16287 20857 16288
rect 3395 15808 3711 15809
rect 3395 15744 3401 15808
rect 3465 15744 3481 15808
rect 3545 15744 3561 15808
rect 3625 15744 3641 15808
rect 3705 15744 3711 15808
rect 3395 15743 3711 15744
rect 8294 15808 8610 15809
rect 8294 15744 8300 15808
rect 8364 15744 8380 15808
rect 8444 15744 8460 15808
rect 8524 15744 8540 15808
rect 8604 15744 8610 15808
rect 8294 15743 8610 15744
rect 13193 15808 13509 15809
rect 13193 15744 13199 15808
rect 13263 15744 13279 15808
rect 13343 15744 13359 15808
rect 13423 15744 13439 15808
rect 13503 15744 13509 15808
rect 13193 15743 13509 15744
rect 18092 15808 18408 15809
rect 18092 15744 18098 15808
rect 18162 15744 18178 15808
rect 18242 15744 18258 15808
rect 18322 15744 18338 15808
rect 18402 15744 18408 15808
rect 18092 15743 18408 15744
rect 19977 15602 20043 15605
rect 21061 15602 21861 15632
rect 19977 15600 21861 15602
rect 19977 15544 19982 15600
rect 20038 15544 21861 15600
rect 19977 15542 21861 15544
rect 19977 15539 20043 15542
rect 21061 15512 21861 15542
rect 5844 15264 6160 15265
rect 5844 15200 5850 15264
rect 5914 15200 5930 15264
rect 5994 15200 6010 15264
rect 6074 15200 6090 15264
rect 6154 15200 6160 15264
rect 5844 15199 6160 15200
rect 10743 15264 11059 15265
rect 10743 15200 10749 15264
rect 10813 15200 10829 15264
rect 10893 15200 10909 15264
rect 10973 15200 10989 15264
rect 11053 15200 11059 15264
rect 10743 15199 11059 15200
rect 15642 15264 15958 15265
rect 15642 15200 15648 15264
rect 15712 15200 15728 15264
rect 15792 15200 15808 15264
rect 15872 15200 15888 15264
rect 15952 15200 15958 15264
rect 15642 15199 15958 15200
rect 20541 15264 20857 15265
rect 20541 15200 20547 15264
rect 20611 15200 20627 15264
rect 20691 15200 20707 15264
rect 20771 15200 20787 15264
rect 20851 15200 20857 15264
rect 20541 15199 20857 15200
rect 3395 14720 3711 14721
rect 3395 14656 3401 14720
rect 3465 14656 3481 14720
rect 3545 14656 3561 14720
rect 3625 14656 3641 14720
rect 3705 14656 3711 14720
rect 3395 14655 3711 14656
rect 8294 14720 8610 14721
rect 8294 14656 8300 14720
rect 8364 14656 8380 14720
rect 8444 14656 8460 14720
rect 8524 14656 8540 14720
rect 8604 14656 8610 14720
rect 8294 14655 8610 14656
rect 13193 14720 13509 14721
rect 13193 14656 13199 14720
rect 13263 14656 13279 14720
rect 13343 14656 13359 14720
rect 13423 14656 13439 14720
rect 13503 14656 13509 14720
rect 13193 14655 13509 14656
rect 18092 14720 18408 14721
rect 18092 14656 18098 14720
rect 18162 14656 18178 14720
rect 18242 14656 18258 14720
rect 18322 14656 18338 14720
rect 18402 14656 18408 14720
rect 18092 14655 18408 14656
rect 5844 14176 6160 14177
rect 5844 14112 5850 14176
rect 5914 14112 5930 14176
rect 5994 14112 6010 14176
rect 6074 14112 6090 14176
rect 6154 14112 6160 14176
rect 5844 14111 6160 14112
rect 10743 14176 11059 14177
rect 10743 14112 10749 14176
rect 10813 14112 10829 14176
rect 10893 14112 10909 14176
rect 10973 14112 10989 14176
rect 11053 14112 11059 14176
rect 10743 14111 11059 14112
rect 15642 14176 15958 14177
rect 15642 14112 15648 14176
rect 15712 14112 15728 14176
rect 15792 14112 15808 14176
rect 15872 14112 15888 14176
rect 15952 14112 15958 14176
rect 15642 14111 15958 14112
rect 20541 14176 20857 14177
rect 20541 14112 20547 14176
rect 20611 14112 20627 14176
rect 20691 14112 20707 14176
rect 20771 14112 20787 14176
rect 20851 14112 20857 14176
rect 20541 14111 20857 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 19977 13834 20043 13837
rect 21061 13834 21861 13864
rect 19977 13832 21861 13834
rect 19977 13776 19982 13832
rect 20038 13776 21861 13832
rect 19977 13774 21861 13776
rect 19977 13771 20043 13774
rect 21061 13744 21861 13774
rect 3395 13632 3711 13633
rect 3395 13568 3401 13632
rect 3465 13568 3481 13632
rect 3545 13568 3561 13632
rect 3625 13568 3641 13632
rect 3705 13568 3711 13632
rect 3395 13567 3711 13568
rect 8294 13632 8610 13633
rect 8294 13568 8300 13632
rect 8364 13568 8380 13632
rect 8444 13568 8460 13632
rect 8524 13568 8540 13632
rect 8604 13568 8610 13632
rect 8294 13567 8610 13568
rect 13193 13632 13509 13633
rect 13193 13568 13199 13632
rect 13263 13568 13279 13632
rect 13343 13568 13359 13632
rect 13423 13568 13439 13632
rect 13503 13568 13509 13632
rect 13193 13567 13509 13568
rect 18092 13632 18408 13633
rect 18092 13568 18098 13632
rect 18162 13568 18178 13632
rect 18242 13568 18258 13632
rect 18322 13568 18338 13632
rect 18402 13568 18408 13632
rect 18092 13567 18408 13568
rect 5844 13088 6160 13089
rect 5844 13024 5850 13088
rect 5914 13024 5930 13088
rect 5994 13024 6010 13088
rect 6074 13024 6090 13088
rect 6154 13024 6160 13088
rect 5844 13023 6160 13024
rect 10743 13088 11059 13089
rect 10743 13024 10749 13088
rect 10813 13024 10829 13088
rect 10893 13024 10909 13088
rect 10973 13024 10989 13088
rect 11053 13024 11059 13088
rect 10743 13023 11059 13024
rect 15642 13088 15958 13089
rect 15642 13024 15648 13088
rect 15712 13024 15728 13088
rect 15792 13024 15808 13088
rect 15872 13024 15888 13088
rect 15952 13024 15958 13088
rect 15642 13023 15958 13024
rect 20541 13088 20857 13089
rect 20541 13024 20547 13088
rect 20611 13024 20627 13088
rect 20691 13024 20707 13088
rect 20771 13024 20787 13088
rect 20851 13024 20857 13088
rect 20541 13023 20857 13024
rect 3395 12544 3711 12545
rect 3395 12480 3401 12544
rect 3465 12480 3481 12544
rect 3545 12480 3561 12544
rect 3625 12480 3641 12544
rect 3705 12480 3711 12544
rect 3395 12479 3711 12480
rect 8294 12544 8610 12545
rect 8294 12480 8300 12544
rect 8364 12480 8380 12544
rect 8444 12480 8460 12544
rect 8524 12480 8540 12544
rect 8604 12480 8610 12544
rect 8294 12479 8610 12480
rect 13193 12544 13509 12545
rect 13193 12480 13199 12544
rect 13263 12480 13279 12544
rect 13343 12480 13359 12544
rect 13423 12480 13439 12544
rect 13503 12480 13509 12544
rect 13193 12479 13509 12480
rect 18092 12544 18408 12545
rect 18092 12480 18098 12544
rect 18162 12480 18178 12544
rect 18242 12480 18258 12544
rect 18322 12480 18338 12544
rect 18402 12480 18408 12544
rect 18092 12479 18408 12480
rect 19977 12338 20043 12341
rect 19977 12336 21466 12338
rect 19977 12280 19982 12336
rect 20038 12280 21466 12336
rect 19977 12278 21466 12280
rect 19977 12275 20043 12278
rect 21406 12096 21466 12278
rect 5844 12000 6160 12001
rect 5844 11936 5850 12000
rect 5914 11936 5930 12000
rect 5994 11936 6010 12000
rect 6074 11936 6090 12000
rect 6154 11936 6160 12000
rect 5844 11935 6160 11936
rect 10743 12000 11059 12001
rect 10743 11936 10749 12000
rect 10813 11936 10829 12000
rect 10893 11936 10909 12000
rect 10973 11936 10989 12000
rect 11053 11936 11059 12000
rect 10743 11935 11059 11936
rect 15642 12000 15958 12001
rect 15642 11936 15648 12000
rect 15712 11936 15728 12000
rect 15792 11936 15808 12000
rect 15872 11936 15888 12000
rect 15952 11936 15958 12000
rect 15642 11935 15958 11936
rect 20541 12000 20857 12001
rect 20541 11936 20547 12000
rect 20611 11936 20627 12000
rect 20691 11936 20707 12000
rect 20771 11936 20787 12000
rect 20851 11936 20857 12000
rect 21061 11976 21861 12096
rect 20541 11935 20857 11936
rect 3395 11456 3711 11457
rect 3395 11392 3401 11456
rect 3465 11392 3481 11456
rect 3545 11392 3561 11456
rect 3625 11392 3641 11456
rect 3705 11392 3711 11456
rect 3395 11391 3711 11392
rect 8294 11456 8610 11457
rect 8294 11392 8300 11456
rect 8364 11392 8380 11456
rect 8444 11392 8460 11456
rect 8524 11392 8540 11456
rect 8604 11392 8610 11456
rect 8294 11391 8610 11392
rect 13193 11456 13509 11457
rect 13193 11392 13199 11456
rect 13263 11392 13279 11456
rect 13343 11392 13359 11456
rect 13423 11392 13439 11456
rect 13503 11392 13509 11456
rect 13193 11391 13509 11392
rect 18092 11456 18408 11457
rect 18092 11392 18098 11456
rect 18162 11392 18178 11456
rect 18242 11392 18258 11456
rect 18322 11392 18338 11456
rect 18402 11392 18408 11456
rect 18092 11391 18408 11392
rect 5844 10912 6160 10913
rect 5844 10848 5850 10912
rect 5914 10848 5930 10912
rect 5994 10848 6010 10912
rect 6074 10848 6090 10912
rect 6154 10848 6160 10912
rect 5844 10847 6160 10848
rect 10743 10912 11059 10913
rect 10743 10848 10749 10912
rect 10813 10848 10829 10912
rect 10893 10848 10909 10912
rect 10973 10848 10989 10912
rect 11053 10848 11059 10912
rect 10743 10847 11059 10848
rect 15642 10912 15958 10913
rect 15642 10848 15648 10912
rect 15712 10848 15728 10912
rect 15792 10848 15808 10912
rect 15872 10848 15888 10912
rect 15952 10848 15958 10912
rect 15642 10847 15958 10848
rect 20541 10912 20857 10913
rect 20541 10848 20547 10912
rect 20611 10848 20627 10912
rect 20691 10848 20707 10912
rect 20771 10848 20787 10912
rect 20851 10848 20857 10912
rect 20541 10847 20857 10848
rect 3395 10368 3711 10369
rect 3395 10304 3401 10368
rect 3465 10304 3481 10368
rect 3545 10304 3561 10368
rect 3625 10304 3641 10368
rect 3705 10304 3711 10368
rect 3395 10303 3711 10304
rect 8294 10368 8610 10369
rect 8294 10304 8300 10368
rect 8364 10304 8380 10368
rect 8444 10304 8460 10368
rect 8524 10304 8540 10368
rect 8604 10304 8610 10368
rect 8294 10303 8610 10304
rect 13193 10368 13509 10369
rect 13193 10304 13199 10368
rect 13263 10304 13279 10368
rect 13343 10304 13359 10368
rect 13423 10304 13439 10368
rect 13503 10304 13509 10368
rect 13193 10303 13509 10304
rect 18092 10368 18408 10369
rect 18092 10304 18098 10368
rect 18162 10304 18178 10368
rect 18242 10304 18258 10368
rect 18322 10304 18338 10368
rect 18402 10304 18408 10368
rect 18092 10303 18408 10304
rect 19977 10298 20043 10301
rect 21061 10298 21861 10328
rect 19977 10296 21861 10298
rect 19977 10240 19982 10296
rect 20038 10240 21861 10296
rect 19977 10238 21861 10240
rect 19977 10235 20043 10238
rect 21061 10208 21861 10238
rect 0 10026 800 10056
rect 1577 10026 1643 10029
rect 0 10024 1643 10026
rect 0 9968 1582 10024
rect 1638 9968 1643 10024
rect 0 9966 1643 9968
rect 0 9936 800 9966
rect 1577 9963 1643 9966
rect 5844 9824 6160 9825
rect 5844 9760 5850 9824
rect 5914 9760 5930 9824
rect 5994 9760 6010 9824
rect 6074 9760 6090 9824
rect 6154 9760 6160 9824
rect 5844 9759 6160 9760
rect 10743 9824 11059 9825
rect 10743 9760 10749 9824
rect 10813 9760 10829 9824
rect 10893 9760 10909 9824
rect 10973 9760 10989 9824
rect 11053 9760 11059 9824
rect 10743 9759 11059 9760
rect 15642 9824 15958 9825
rect 15642 9760 15648 9824
rect 15712 9760 15728 9824
rect 15792 9760 15808 9824
rect 15872 9760 15888 9824
rect 15952 9760 15958 9824
rect 15642 9759 15958 9760
rect 20541 9824 20857 9825
rect 20541 9760 20547 9824
rect 20611 9760 20627 9824
rect 20691 9760 20707 9824
rect 20771 9760 20787 9824
rect 20851 9760 20857 9824
rect 20541 9759 20857 9760
rect 3395 9280 3711 9281
rect 3395 9216 3401 9280
rect 3465 9216 3481 9280
rect 3545 9216 3561 9280
rect 3625 9216 3641 9280
rect 3705 9216 3711 9280
rect 3395 9215 3711 9216
rect 8294 9280 8610 9281
rect 8294 9216 8300 9280
rect 8364 9216 8380 9280
rect 8444 9216 8460 9280
rect 8524 9216 8540 9280
rect 8604 9216 8610 9280
rect 8294 9215 8610 9216
rect 13193 9280 13509 9281
rect 13193 9216 13199 9280
rect 13263 9216 13279 9280
rect 13343 9216 13359 9280
rect 13423 9216 13439 9280
rect 13503 9216 13509 9280
rect 13193 9215 13509 9216
rect 18092 9280 18408 9281
rect 18092 9216 18098 9280
rect 18162 9216 18178 9280
rect 18242 9216 18258 9280
rect 18322 9216 18338 9280
rect 18402 9216 18408 9280
rect 18092 9215 18408 9216
rect 5844 8736 6160 8737
rect 5844 8672 5850 8736
rect 5914 8672 5930 8736
rect 5994 8672 6010 8736
rect 6074 8672 6090 8736
rect 6154 8672 6160 8736
rect 5844 8671 6160 8672
rect 10743 8736 11059 8737
rect 10743 8672 10749 8736
rect 10813 8672 10829 8736
rect 10893 8672 10909 8736
rect 10973 8672 10989 8736
rect 11053 8672 11059 8736
rect 10743 8671 11059 8672
rect 15642 8736 15958 8737
rect 15642 8672 15648 8736
rect 15712 8672 15728 8736
rect 15792 8672 15808 8736
rect 15872 8672 15888 8736
rect 15952 8672 15958 8736
rect 15642 8671 15958 8672
rect 20541 8736 20857 8737
rect 20541 8672 20547 8736
rect 20611 8672 20627 8736
rect 20691 8672 20707 8736
rect 20771 8672 20787 8736
rect 20851 8672 20857 8736
rect 20541 8671 20857 8672
rect 19977 8530 20043 8533
rect 21061 8530 21861 8560
rect 19977 8528 21861 8530
rect 19977 8472 19982 8528
rect 20038 8472 21861 8528
rect 19977 8470 21861 8472
rect 19977 8467 20043 8470
rect 21061 8440 21861 8470
rect 3395 8192 3711 8193
rect 3395 8128 3401 8192
rect 3465 8128 3481 8192
rect 3545 8128 3561 8192
rect 3625 8128 3641 8192
rect 3705 8128 3711 8192
rect 3395 8127 3711 8128
rect 8294 8192 8610 8193
rect 8294 8128 8300 8192
rect 8364 8128 8380 8192
rect 8444 8128 8460 8192
rect 8524 8128 8540 8192
rect 8604 8128 8610 8192
rect 8294 8127 8610 8128
rect 13193 8192 13509 8193
rect 13193 8128 13199 8192
rect 13263 8128 13279 8192
rect 13343 8128 13359 8192
rect 13423 8128 13439 8192
rect 13503 8128 13509 8192
rect 13193 8127 13509 8128
rect 18092 8192 18408 8193
rect 18092 8128 18098 8192
rect 18162 8128 18178 8192
rect 18242 8128 18258 8192
rect 18322 8128 18338 8192
rect 18402 8128 18408 8192
rect 18092 8127 18408 8128
rect 5844 7648 6160 7649
rect 5844 7584 5850 7648
rect 5914 7584 5930 7648
rect 5994 7584 6010 7648
rect 6074 7584 6090 7648
rect 6154 7584 6160 7648
rect 5844 7583 6160 7584
rect 10743 7648 11059 7649
rect 10743 7584 10749 7648
rect 10813 7584 10829 7648
rect 10893 7584 10909 7648
rect 10973 7584 10989 7648
rect 11053 7584 11059 7648
rect 10743 7583 11059 7584
rect 15642 7648 15958 7649
rect 15642 7584 15648 7648
rect 15712 7584 15728 7648
rect 15792 7584 15808 7648
rect 15872 7584 15888 7648
rect 15952 7584 15958 7648
rect 15642 7583 15958 7584
rect 20541 7648 20857 7649
rect 20541 7584 20547 7648
rect 20611 7584 20627 7648
rect 20691 7584 20707 7648
rect 20771 7584 20787 7648
rect 20851 7584 20857 7648
rect 20541 7583 20857 7584
rect 3395 7104 3711 7105
rect 3395 7040 3401 7104
rect 3465 7040 3481 7104
rect 3545 7040 3561 7104
rect 3625 7040 3641 7104
rect 3705 7040 3711 7104
rect 3395 7039 3711 7040
rect 8294 7104 8610 7105
rect 8294 7040 8300 7104
rect 8364 7040 8380 7104
rect 8444 7040 8460 7104
rect 8524 7040 8540 7104
rect 8604 7040 8610 7104
rect 8294 7039 8610 7040
rect 13193 7104 13509 7105
rect 13193 7040 13199 7104
rect 13263 7040 13279 7104
rect 13343 7040 13359 7104
rect 13423 7040 13439 7104
rect 13503 7040 13509 7104
rect 13193 7039 13509 7040
rect 18092 7104 18408 7105
rect 18092 7040 18098 7104
rect 18162 7040 18178 7104
rect 18242 7040 18258 7104
rect 18322 7040 18338 7104
rect 18402 7040 18408 7104
rect 18092 7039 18408 7040
rect 19977 6762 20043 6765
rect 21061 6762 21861 6792
rect 19977 6760 21861 6762
rect 19977 6704 19982 6760
rect 20038 6704 21861 6760
rect 19977 6702 21861 6704
rect 19977 6699 20043 6702
rect 21061 6672 21861 6702
rect 5844 6560 6160 6561
rect 5844 6496 5850 6560
rect 5914 6496 5930 6560
rect 5994 6496 6010 6560
rect 6074 6496 6090 6560
rect 6154 6496 6160 6560
rect 5844 6495 6160 6496
rect 10743 6560 11059 6561
rect 10743 6496 10749 6560
rect 10813 6496 10829 6560
rect 10893 6496 10909 6560
rect 10973 6496 10989 6560
rect 11053 6496 11059 6560
rect 10743 6495 11059 6496
rect 15642 6560 15958 6561
rect 15642 6496 15648 6560
rect 15712 6496 15728 6560
rect 15792 6496 15808 6560
rect 15872 6496 15888 6560
rect 15952 6496 15958 6560
rect 15642 6495 15958 6496
rect 20541 6560 20857 6561
rect 20541 6496 20547 6560
rect 20611 6496 20627 6560
rect 20691 6496 20707 6560
rect 20771 6496 20787 6560
rect 20851 6496 20857 6560
rect 20541 6495 20857 6496
rect 0 6100 800 6112
rect 0 6017 3700 6100
rect 0 6016 3711 6017
rect 0 6000 3401 6016
rect 0 5992 800 6000
rect 3395 5952 3401 6000
rect 3465 5952 3481 6016
rect 3545 5952 3561 6016
rect 3625 5952 3641 6016
rect 3705 5952 3711 6016
rect 3395 5951 3711 5952
rect 8294 6016 8610 6017
rect 8294 5952 8300 6016
rect 8364 5952 8380 6016
rect 8444 5952 8460 6016
rect 8524 5952 8540 6016
rect 8604 5952 8610 6016
rect 8294 5951 8610 5952
rect 13193 6016 13509 6017
rect 13193 5952 13199 6016
rect 13263 5952 13279 6016
rect 13343 5952 13359 6016
rect 13423 5952 13439 6016
rect 13503 5952 13509 6016
rect 13193 5951 13509 5952
rect 18092 6016 18408 6017
rect 18092 5952 18098 6016
rect 18162 5952 18178 6016
rect 18242 5952 18258 6016
rect 18322 5952 18338 6016
rect 18402 5952 18408 6016
rect 18092 5951 18408 5952
rect 5844 5472 6160 5473
rect 5844 5408 5850 5472
rect 5914 5408 5930 5472
rect 5994 5408 6010 5472
rect 6074 5408 6090 5472
rect 6154 5408 6160 5472
rect 5844 5407 6160 5408
rect 10743 5472 11059 5473
rect 10743 5408 10749 5472
rect 10813 5408 10829 5472
rect 10893 5408 10909 5472
rect 10973 5408 10989 5472
rect 11053 5408 11059 5472
rect 10743 5407 11059 5408
rect 15642 5472 15958 5473
rect 15642 5408 15648 5472
rect 15712 5408 15728 5472
rect 15792 5408 15808 5472
rect 15872 5408 15888 5472
rect 15952 5408 15958 5472
rect 15642 5407 15958 5408
rect 20541 5472 20857 5473
rect 20541 5408 20547 5472
rect 20611 5408 20627 5472
rect 20691 5408 20707 5472
rect 20771 5408 20787 5472
rect 20851 5408 20857 5472
rect 20541 5407 20857 5408
rect 20069 4994 20135 4997
rect 21061 4994 21861 5024
rect 20069 4992 21861 4994
rect 20069 4936 20074 4992
rect 20130 4936 21861 4992
rect 20069 4934 21861 4936
rect 20069 4931 20135 4934
rect 3395 4928 3711 4929
rect 3395 4864 3401 4928
rect 3465 4864 3481 4928
rect 3545 4864 3561 4928
rect 3625 4864 3641 4928
rect 3705 4864 3711 4928
rect 3395 4863 3711 4864
rect 8294 4928 8610 4929
rect 8294 4864 8300 4928
rect 8364 4864 8380 4928
rect 8444 4864 8460 4928
rect 8524 4864 8540 4928
rect 8604 4864 8610 4928
rect 8294 4863 8610 4864
rect 13193 4928 13509 4929
rect 13193 4864 13199 4928
rect 13263 4864 13279 4928
rect 13343 4864 13359 4928
rect 13423 4864 13439 4928
rect 13503 4864 13509 4928
rect 13193 4863 13509 4864
rect 18092 4928 18408 4929
rect 18092 4864 18098 4928
rect 18162 4864 18178 4928
rect 18242 4864 18258 4928
rect 18322 4864 18338 4928
rect 18402 4864 18408 4928
rect 21061 4904 21861 4934
rect 18092 4863 18408 4864
rect 5844 4384 6160 4385
rect 5844 4320 5850 4384
rect 5914 4320 5930 4384
rect 5994 4320 6010 4384
rect 6074 4320 6090 4384
rect 6154 4320 6160 4384
rect 5844 4319 6160 4320
rect 10743 4384 11059 4385
rect 10743 4320 10749 4384
rect 10813 4320 10829 4384
rect 10893 4320 10909 4384
rect 10973 4320 10989 4384
rect 11053 4320 11059 4384
rect 10743 4319 11059 4320
rect 15642 4384 15958 4385
rect 15642 4320 15648 4384
rect 15712 4320 15728 4384
rect 15792 4320 15808 4384
rect 15872 4320 15888 4384
rect 15952 4320 15958 4384
rect 15642 4319 15958 4320
rect 20541 4384 20857 4385
rect 20541 4320 20547 4384
rect 20611 4320 20627 4384
rect 20691 4320 20707 4384
rect 20771 4320 20787 4384
rect 20851 4320 20857 4384
rect 20541 4319 20857 4320
rect 3395 3840 3711 3841
rect 3395 3776 3401 3840
rect 3465 3776 3481 3840
rect 3545 3776 3561 3840
rect 3625 3776 3641 3840
rect 3705 3776 3711 3840
rect 3395 3775 3711 3776
rect 8294 3840 8610 3841
rect 8294 3776 8300 3840
rect 8364 3776 8380 3840
rect 8444 3776 8460 3840
rect 8524 3776 8540 3840
rect 8604 3776 8610 3840
rect 8294 3775 8610 3776
rect 13193 3840 13509 3841
rect 13193 3776 13199 3840
rect 13263 3776 13279 3840
rect 13343 3776 13359 3840
rect 13423 3776 13439 3840
rect 13503 3776 13509 3840
rect 13193 3775 13509 3776
rect 18092 3840 18408 3841
rect 18092 3776 18098 3840
rect 18162 3776 18178 3840
rect 18242 3776 18258 3840
rect 18322 3776 18338 3840
rect 18402 3776 18408 3840
rect 18092 3775 18408 3776
rect 20069 3498 20135 3501
rect 21214 3498 21220 3500
rect 20069 3496 21220 3498
rect 20069 3440 20074 3496
rect 20130 3440 21220 3496
rect 20069 3438 21220 3440
rect 20069 3435 20135 3438
rect 21214 3436 21220 3438
rect 21284 3436 21290 3500
rect 5844 3296 6160 3297
rect 5844 3232 5850 3296
rect 5914 3232 5930 3296
rect 5994 3232 6010 3296
rect 6074 3232 6090 3296
rect 6154 3232 6160 3296
rect 5844 3231 6160 3232
rect 10743 3296 11059 3297
rect 10743 3232 10749 3296
rect 10813 3232 10829 3296
rect 10893 3232 10909 3296
rect 10973 3232 10989 3296
rect 11053 3232 11059 3296
rect 10743 3231 11059 3232
rect 15642 3296 15958 3297
rect 15642 3232 15648 3296
rect 15712 3232 15728 3296
rect 15792 3232 15808 3296
rect 15872 3232 15888 3296
rect 15952 3232 15958 3296
rect 15642 3231 15958 3232
rect 20541 3296 20857 3297
rect 20541 3232 20547 3296
rect 20611 3232 20627 3296
rect 20691 3232 20707 3296
rect 20771 3232 20787 3296
rect 20851 3232 20857 3296
rect 20541 3231 20857 3232
rect 21061 3228 21861 3256
rect 21061 3164 21220 3228
rect 21284 3164 21861 3228
rect 21061 3136 21861 3164
rect 3395 2752 3711 2753
rect 3395 2688 3401 2752
rect 3465 2688 3481 2752
rect 3545 2688 3561 2752
rect 3625 2688 3641 2752
rect 3705 2688 3711 2752
rect 3395 2687 3711 2688
rect 8294 2752 8610 2753
rect 8294 2688 8300 2752
rect 8364 2688 8380 2752
rect 8444 2688 8460 2752
rect 8524 2688 8540 2752
rect 8604 2688 8610 2752
rect 8294 2687 8610 2688
rect 13193 2752 13509 2753
rect 13193 2688 13199 2752
rect 13263 2688 13279 2752
rect 13343 2688 13359 2752
rect 13423 2688 13439 2752
rect 13503 2688 13509 2752
rect 13193 2687 13509 2688
rect 18092 2752 18408 2753
rect 18092 2688 18098 2752
rect 18162 2688 18178 2752
rect 18242 2688 18258 2752
rect 18322 2688 18338 2752
rect 18402 2688 18408 2752
rect 18092 2687 18408 2688
rect 5844 2208 6160 2209
rect 0 2138 800 2168
rect 5844 2144 5850 2208
rect 5914 2144 5930 2208
rect 5994 2144 6010 2208
rect 6074 2144 6090 2208
rect 6154 2144 6160 2208
rect 5844 2143 6160 2144
rect 10743 2208 11059 2209
rect 10743 2144 10749 2208
rect 10813 2144 10829 2208
rect 10893 2144 10909 2208
rect 10973 2144 10989 2208
rect 11053 2144 11059 2208
rect 10743 2143 11059 2144
rect 15642 2208 15958 2209
rect 15642 2144 15648 2208
rect 15712 2144 15728 2208
rect 15792 2144 15808 2208
rect 15872 2144 15888 2208
rect 15952 2144 15958 2208
rect 15642 2143 15958 2144
rect 20541 2208 20857 2209
rect 20541 2144 20547 2208
rect 20611 2144 20627 2208
rect 20691 2144 20707 2208
rect 20771 2144 20787 2208
rect 20851 2144 20857 2208
rect 20541 2143 20857 2144
rect 1761 2138 1827 2141
rect 0 2136 1827 2138
rect 0 2080 1766 2136
rect 1822 2080 1827 2136
rect 0 2078 1827 2080
rect 0 2048 800 2078
rect 1761 2075 1827 2078
rect 19149 1458 19215 1461
rect 21061 1458 21861 1488
rect 19149 1456 21861 1458
rect 19149 1400 19154 1456
rect 19210 1400 21861 1456
rect 19149 1398 21861 1400
rect 19149 1395 19215 1398
rect 21061 1368 21861 1398
<< via3 >>
rect 5850 21788 5914 21792
rect 5850 21732 5854 21788
rect 5854 21732 5910 21788
rect 5910 21732 5914 21788
rect 5850 21728 5914 21732
rect 5930 21788 5994 21792
rect 5930 21732 5934 21788
rect 5934 21732 5990 21788
rect 5990 21732 5994 21788
rect 5930 21728 5994 21732
rect 6010 21788 6074 21792
rect 6010 21732 6014 21788
rect 6014 21732 6070 21788
rect 6070 21732 6074 21788
rect 6010 21728 6074 21732
rect 6090 21788 6154 21792
rect 6090 21732 6094 21788
rect 6094 21732 6150 21788
rect 6150 21732 6154 21788
rect 6090 21728 6154 21732
rect 10749 21788 10813 21792
rect 10749 21732 10753 21788
rect 10753 21732 10809 21788
rect 10809 21732 10813 21788
rect 10749 21728 10813 21732
rect 10829 21788 10893 21792
rect 10829 21732 10833 21788
rect 10833 21732 10889 21788
rect 10889 21732 10893 21788
rect 10829 21728 10893 21732
rect 10909 21788 10973 21792
rect 10909 21732 10913 21788
rect 10913 21732 10969 21788
rect 10969 21732 10973 21788
rect 10909 21728 10973 21732
rect 10989 21788 11053 21792
rect 10989 21732 10993 21788
rect 10993 21732 11049 21788
rect 11049 21732 11053 21788
rect 10989 21728 11053 21732
rect 15648 21788 15712 21792
rect 15648 21732 15652 21788
rect 15652 21732 15708 21788
rect 15708 21732 15712 21788
rect 15648 21728 15712 21732
rect 15728 21788 15792 21792
rect 15728 21732 15732 21788
rect 15732 21732 15788 21788
rect 15788 21732 15792 21788
rect 15728 21728 15792 21732
rect 15808 21788 15872 21792
rect 15808 21732 15812 21788
rect 15812 21732 15868 21788
rect 15868 21732 15872 21788
rect 15808 21728 15872 21732
rect 15888 21788 15952 21792
rect 15888 21732 15892 21788
rect 15892 21732 15948 21788
rect 15948 21732 15952 21788
rect 15888 21728 15952 21732
rect 20547 21788 20611 21792
rect 20547 21732 20551 21788
rect 20551 21732 20607 21788
rect 20607 21732 20611 21788
rect 20547 21728 20611 21732
rect 20627 21788 20691 21792
rect 20627 21732 20631 21788
rect 20631 21732 20687 21788
rect 20687 21732 20691 21788
rect 20627 21728 20691 21732
rect 20707 21788 20771 21792
rect 20707 21732 20711 21788
rect 20711 21732 20767 21788
rect 20767 21732 20771 21788
rect 20707 21728 20771 21732
rect 20787 21788 20851 21792
rect 20787 21732 20791 21788
rect 20791 21732 20847 21788
rect 20847 21732 20851 21788
rect 20787 21728 20851 21732
rect 3401 21244 3465 21248
rect 3401 21188 3405 21244
rect 3405 21188 3461 21244
rect 3461 21188 3465 21244
rect 3401 21184 3465 21188
rect 3481 21244 3545 21248
rect 3481 21188 3485 21244
rect 3485 21188 3541 21244
rect 3541 21188 3545 21244
rect 3481 21184 3545 21188
rect 3561 21244 3625 21248
rect 3561 21188 3565 21244
rect 3565 21188 3621 21244
rect 3621 21188 3625 21244
rect 3561 21184 3625 21188
rect 3641 21244 3705 21248
rect 3641 21188 3645 21244
rect 3645 21188 3701 21244
rect 3701 21188 3705 21244
rect 3641 21184 3705 21188
rect 8300 21244 8364 21248
rect 8300 21188 8304 21244
rect 8304 21188 8360 21244
rect 8360 21188 8364 21244
rect 8300 21184 8364 21188
rect 8380 21244 8444 21248
rect 8380 21188 8384 21244
rect 8384 21188 8440 21244
rect 8440 21188 8444 21244
rect 8380 21184 8444 21188
rect 8460 21244 8524 21248
rect 8460 21188 8464 21244
rect 8464 21188 8520 21244
rect 8520 21188 8524 21244
rect 8460 21184 8524 21188
rect 8540 21244 8604 21248
rect 8540 21188 8544 21244
rect 8544 21188 8600 21244
rect 8600 21188 8604 21244
rect 8540 21184 8604 21188
rect 13199 21244 13263 21248
rect 13199 21188 13203 21244
rect 13203 21188 13259 21244
rect 13259 21188 13263 21244
rect 13199 21184 13263 21188
rect 13279 21244 13343 21248
rect 13279 21188 13283 21244
rect 13283 21188 13339 21244
rect 13339 21188 13343 21244
rect 13279 21184 13343 21188
rect 13359 21244 13423 21248
rect 13359 21188 13363 21244
rect 13363 21188 13419 21244
rect 13419 21188 13423 21244
rect 13359 21184 13423 21188
rect 13439 21244 13503 21248
rect 13439 21188 13443 21244
rect 13443 21188 13499 21244
rect 13499 21188 13503 21244
rect 13439 21184 13503 21188
rect 18098 21244 18162 21248
rect 18098 21188 18102 21244
rect 18102 21188 18158 21244
rect 18158 21188 18162 21244
rect 18098 21184 18162 21188
rect 18178 21244 18242 21248
rect 18178 21188 18182 21244
rect 18182 21188 18238 21244
rect 18238 21188 18242 21244
rect 18178 21184 18242 21188
rect 18258 21244 18322 21248
rect 18258 21188 18262 21244
rect 18262 21188 18318 21244
rect 18318 21188 18322 21244
rect 18258 21184 18322 21188
rect 18338 21244 18402 21248
rect 18338 21188 18342 21244
rect 18342 21188 18398 21244
rect 18398 21188 18402 21244
rect 18338 21184 18402 21188
rect 5850 20700 5914 20704
rect 5850 20644 5854 20700
rect 5854 20644 5910 20700
rect 5910 20644 5914 20700
rect 5850 20640 5914 20644
rect 5930 20700 5994 20704
rect 5930 20644 5934 20700
rect 5934 20644 5990 20700
rect 5990 20644 5994 20700
rect 5930 20640 5994 20644
rect 6010 20700 6074 20704
rect 6010 20644 6014 20700
rect 6014 20644 6070 20700
rect 6070 20644 6074 20700
rect 6010 20640 6074 20644
rect 6090 20700 6154 20704
rect 6090 20644 6094 20700
rect 6094 20644 6150 20700
rect 6150 20644 6154 20700
rect 6090 20640 6154 20644
rect 10749 20700 10813 20704
rect 10749 20644 10753 20700
rect 10753 20644 10809 20700
rect 10809 20644 10813 20700
rect 10749 20640 10813 20644
rect 10829 20700 10893 20704
rect 10829 20644 10833 20700
rect 10833 20644 10889 20700
rect 10889 20644 10893 20700
rect 10829 20640 10893 20644
rect 10909 20700 10973 20704
rect 10909 20644 10913 20700
rect 10913 20644 10969 20700
rect 10969 20644 10973 20700
rect 10909 20640 10973 20644
rect 10989 20700 11053 20704
rect 10989 20644 10993 20700
rect 10993 20644 11049 20700
rect 11049 20644 11053 20700
rect 10989 20640 11053 20644
rect 15648 20700 15712 20704
rect 15648 20644 15652 20700
rect 15652 20644 15708 20700
rect 15708 20644 15712 20700
rect 15648 20640 15712 20644
rect 15728 20700 15792 20704
rect 15728 20644 15732 20700
rect 15732 20644 15788 20700
rect 15788 20644 15792 20700
rect 15728 20640 15792 20644
rect 15808 20700 15872 20704
rect 15808 20644 15812 20700
rect 15812 20644 15868 20700
rect 15868 20644 15872 20700
rect 15808 20640 15872 20644
rect 15888 20700 15952 20704
rect 15888 20644 15892 20700
rect 15892 20644 15948 20700
rect 15948 20644 15952 20700
rect 15888 20640 15952 20644
rect 20547 20700 20611 20704
rect 20547 20644 20551 20700
rect 20551 20644 20607 20700
rect 20607 20644 20611 20700
rect 20547 20640 20611 20644
rect 20627 20700 20691 20704
rect 20627 20644 20631 20700
rect 20631 20644 20687 20700
rect 20687 20644 20691 20700
rect 20627 20640 20691 20644
rect 20707 20700 20771 20704
rect 20707 20644 20711 20700
rect 20711 20644 20767 20700
rect 20767 20644 20771 20700
rect 20707 20640 20771 20644
rect 20787 20700 20851 20704
rect 20787 20644 20791 20700
rect 20791 20644 20847 20700
rect 20847 20644 20851 20700
rect 20787 20640 20851 20644
rect 3401 20156 3465 20160
rect 3401 20100 3405 20156
rect 3405 20100 3461 20156
rect 3461 20100 3465 20156
rect 3401 20096 3465 20100
rect 3481 20156 3545 20160
rect 3481 20100 3485 20156
rect 3485 20100 3541 20156
rect 3541 20100 3545 20156
rect 3481 20096 3545 20100
rect 3561 20156 3625 20160
rect 3561 20100 3565 20156
rect 3565 20100 3621 20156
rect 3621 20100 3625 20156
rect 3561 20096 3625 20100
rect 3641 20156 3705 20160
rect 3641 20100 3645 20156
rect 3645 20100 3701 20156
rect 3701 20100 3705 20156
rect 3641 20096 3705 20100
rect 8300 20156 8364 20160
rect 8300 20100 8304 20156
rect 8304 20100 8360 20156
rect 8360 20100 8364 20156
rect 8300 20096 8364 20100
rect 8380 20156 8444 20160
rect 8380 20100 8384 20156
rect 8384 20100 8440 20156
rect 8440 20100 8444 20156
rect 8380 20096 8444 20100
rect 8460 20156 8524 20160
rect 8460 20100 8464 20156
rect 8464 20100 8520 20156
rect 8520 20100 8524 20156
rect 8460 20096 8524 20100
rect 8540 20156 8604 20160
rect 8540 20100 8544 20156
rect 8544 20100 8600 20156
rect 8600 20100 8604 20156
rect 8540 20096 8604 20100
rect 13199 20156 13263 20160
rect 13199 20100 13203 20156
rect 13203 20100 13259 20156
rect 13259 20100 13263 20156
rect 13199 20096 13263 20100
rect 13279 20156 13343 20160
rect 13279 20100 13283 20156
rect 13283 20100 13339 20156
rect 13339 20100 13343 20156
rect 13279 20096 13343 20100
rect 13359 20156 13423 20160
rect 13359 20100 13363 20156
rect 13363 20100 13419 20156
rect 13419 20100 13423 20156
rect 13359 20096 13423 20100
rect 13439 20156 13503 20160
rect 13439 20100 13443 20156
rect 13443 20100 13499 20156
rect 13499 20100 13503 20156
rect 13439 20096 13503 20100
rect 18098 20156 18162 20160
rect 18098 20100 18102 20156
rect 18102 20100 18158 20156
rect 18158 20100 18162 20156
rect 18098 20096 18162 20100
rect 18178 20156 18242 20160
rect 18178 20100 18182 20156
rect 18182 20100 18238 20156
rect 18238 20100 18242 20156
rect 18178 20096 18242 20100
rect 18258 20156 18322 20160
rect 18258 20100 18262 20156
rect 18262 20100 18318 20156
rect 18318 20100 18322 20156
rect 18258 20096 18322 20100
rect 18338 20156 18402 20160
rect 18338 20100 18342 20156
rect 18342 20100 18398 20156
rect 18398 20100 18402 20156
rect 18338 20096 18402 20100
rect 5850 19612 5914 19616
rect 5850 19556 5854 19612
rect 5854 19556 5910 19612
rect 5910 19556 5914 19612
rect 5850 19552 5914 19556
rect 5930 19612 5994 19616
rect 5930 19556 5934 19612
rect 5934 19556 5990 19612
rect 5990 19556 5994 19612
rect 5930 19552 5994 19556
rect 6010 19612 6074 19616
rect 6010 19556 6014 19612
rect 6014 19556 6070 19612
rect 6070 19556 6074 19612
rect 6010 19552 6074 19556
rect 6090 19612 6154 19616
rect 6090 19556 6094 19612
rect 6094 19556 6150 19612
rect 6150 19556 6154 19612
rect 6090 19552 6154 19556
rect 10749 19612 10813 19616
rect 10749 19556 10753 19612
rect 10753 19556 10809 19612
rect 10809 19556 10813 19612
rect 10749 19552 10813 19556
rect 10829 19612 10893 19616
rect 10829 19556 10833 19612
rect 10833 19556 10889 19612
rect 10889 19556 10893 19612
rect 10829 19552 10893 19556
rect 10909 19612 10973 19616
rect 10909 19556 10913 19612
rect 10913 19556 10969 19612
rect 10969 19556 10973 19612
rect 10909 19552 10973 19556
rect 10989 19612 11053 19616
rect 10989 19556 10993 19612
rect 10993 19556 11049 19612
rect 11049 19556 11053 19612
rect 10989 19552 11053 19556
rect 15648 19612 15712 19616
rect 15648 19556 15652 19612
rect 15652 19556 15708 19612
rect 15708 19556 15712 19612
rect 15648 19552 15712 19556
rect 15728 19612 15792 19616
rect 15728 19556 15732 19612
rect 15732 19556 15788 19612
rect 15788 19556 15792 19612
rect 15728 19552 15792 19556
rect 15808 19612 15872 19616
rect 15808 19556 15812 19612
rect 15812 19556 15868 19612
rect 15868 19556 15872 19612
rect 15808 19552 15872 19556
rect 15888 19612 15952 19616
rect 15888 19556 15892 19612
rect 15892 19556 15948 19612
rect 15948 19556 15952 19612
rect 15888 19552 15952 19556
rect 20547 19612 20611 19616
rect 20547 19556 20551 19612
rect 20551 19556 20607 19612
rect 20607 19556 20611 19612
rect 20547 19552 20611 19556
rect 20627 19612 20691 19616
rect 20627 19556 20631 19612
rect 20631 19556 20687 19612
rect 20687 19556 20691 19612
rect 20627 19552 20691 19556
rect 20707 19612 20771 19616
rect 20707 19556 20711 19612
rect 20711 19556 20767 19612
rect 20767 19556 20771 19612
rect 20707 19552 20771 19556
rect 20787 19612 20851 19616
rect 20787 19556 20791 19612
rect 20791 19556 20847 19612
rect 20847 19556 20851 19612
rect 20787 19552 20851 19556
rect 3401 19068 3465 19072
rect 3401 19012 3405 19068
rect 3405 19012 3461 19068
rect 3461 19012 3465 19068
rect 3401 19008 3465 19012
rect 3481 19068 3545 19072
rect 3481 19012 3485 19068
rect 3485 19012 3541 19068
rect 3541 19012 3545 19068
rect 3481 19008 3545 19012
rect 3561 19068 3625 19072
rect 3561 19012 3565 19068
rect 3565 19012 3621 19068
rect 3621 19012 3625 19068
rect 3561 19008 3625 19012
rect 3641 19068 3705 19072
rect 3641 19012 3645 19068
rect 3645 19012 3701 19068
rect 3701 19012 3705 19068
rect 3641 19008 3705 19012
rect 8300 19068 8364 19072
rect 8300 19012 8304 19068
rect 8304 19012 8360 19068
rect 8360 19012 8364 19068
rect 8300 19008 8364 19012
rect 8380 19068 8444 19072
rect 8380 19012 8384 19068
rect 8384 19012 8440 19068
rect 8440 19012 8444 19068
rect 8380 19008 8444 19012
rect 8460 19068 8524 19072
rect 8460 19012 8464 19068
rect 8464 19012 8520 19068
rect 8520 19012 8524 19068
rect 8460 19008 8524 19012
rect 8540 19068 8604 19072
rect 8540 19012 8544 19068
rect 8544 19012 8600 19068
rect 8600 19012 8604 19068
rect 8540 19008 8604 19012
rect 13199 19068 13263 19072
rect 13199 19012 13203 19068
rect 13203 19012 13259 19068
rect 13259 19012 13263 19068
rect 13199 19008 13263 19012
rect 13279 19068 13343 19072
rect 13279 19012 13283 19068
rect 13283 19012 13339 19068
rect 13339 19012 13343 19068
rect 13279 19008 13343 19012
rect 13359 19068 13423 19072
rect 13359 19012 13363 19068
rect 13363 19012 13419 19068
rect 13419 19012 13423 19068
rect 13359 19008 13423 19012
rect 13439 19068 13503 19072
rect 13439 19012 13443 19068
rect 13443 19012 13499 19068
rect 13499 19012 13503 19068
rect 13439 19008 13503 19012
rect 18098 19068 18162 19072
rect 18098 19012 18102 19068
rect 18102 19012 18158 19068
rect 18158 19012 18162 19068
rect 18098 19008 18162 19012
rect 18178 19068 18242 19072
rect 18178 19012 18182 19068
rect 18182 19012 18238 19068
rect 18238 19012 18242 19068
rect 18178 19008 18242 19012
rect 18258 19068 18322 19072
rect 18258 19012 18262 19068
rect 18262 19012 18318 19068
rect 18318 19012 18322 19068
rect 18258 19008 18322 19012
rect 18338 19068 18402 19072
rect 18338 19012 18342 19068
rect 18342 19012 18398 19068
rect 18398 19012 18402 19068
rect 18338 19008 18402 19012
rect 5850 18524 5914 18528
rect 5850 18468 5854 18524
rect 5854 18468 5910 18524
rect 5910 18468 5914 18524
rect 5850 18464 5914 18468
rect 5930 18524 5994 18528
rect 5930 18468 5934 18524
rect 5934 18468 5990 18524
rect 5990 18468 5994 18524
rect 5930 18464 5994 18468
rect 6010 18524 6074 18528
rect 6010 18468 6014 18524
rect 6014 18468 6070 18524
rect 6070 18468 6074 18524
rect 6010 18464 6074 18468
rect 6090 18524 6154 18528
rect 6090 18468 6094 18524
rect 6094 18468 6150 18524
rect 6150 18468 6154 18524
rect 6090 18464 6154 18468
rect 10749 18524 10813 18528
rect 10749 18468 10753 18524
rect 10753 18468 10809 18524
rect 10809 18468 10813 18524
rect 10749 18464 10813 18468
rect 10829 18524 10893 18528
rect 10829 18468 10833 18524
rect 10833 18468 10889 18524
rect 10889 18468 10893 18524
rect 10829 18464 10893 18468
rect 10909 18524 10973 18528
rect 10909 18468 10913 18524
rect 10913 18468 10969 18524
rect 10969 18468 10973 18524
rect 10909 18464 10973 18468
rect 10989 18524 11053 18528
rect 10989 18468 10993 18524
rect 10993 18468 11049 18524
rect 11049 18468 11053 18524
rect 10989 18464 11053 18468
rect 15648 18524 15712 18528
rect 15648 18468 15652 18524
rect 15652 18468 15708 18524
rect 15708 18468 15712 18524
rect 15648 18464 15712 18468
rect 15728 18524 15792 18528
rect 15728 18468 15732 18524
rect 15732 18468 15788 18524
rect 15788 18468 15792 18524
rect 15728 18464 15792 18468
rect 15808 18524 15872 18528
rect 15808 18468 15812 18524
rect 15812 18468 15868 18524
rect 15868 18468 15872 18524
rect 15808 18464 15872 18468
rect 15888 18524 15952 18528
rect 15888 18468 15892 18524
rect 15892 18468 15948 18524
rect 15948 18468 15952 18524
rect 15888 18464 15952 18468
rect 20547 18524 20611 18528
rect 20547 18468 20551 18524
rect 20551 18468 20607 18524
rect 20607 18468 20611 18524
rect 20547 18464 20611 18468
rect 20627 18524 20691 18528
rect 20627 18468 20631 18524
rect 20631 18468 20687 18524
rect 20687 18468 20691 18524
rect 20627 18464 20691 18468
rect 20707 18524 20771 18528
rect 20707 18468 20711 18524
rect 20711 18468 20767 18524
rect 20767 18468 20771 18524
rect 20707 18464 20771 18468
rect 20787 18524 20851 18528
rect 20787 18468 20791 18524
rect 20791 18468 20847 18524
rect 20847 18468 20851 18524
rect 20787 18464 20851 18468
rect 3401 17980 3465 17984
rect 3401 17924 3405 17980
rect 3405 17924 3461 17980
rect 3461 17924 3465 17980
rect 3401 17920 3465 17924
rect 3481 17980 3545 17984
rect 3481 17924 3485 17980
rect 3485 17924 3541 17980
rect 3541 17924 3545 17980
rect 3481 17920 3545 17924
rect 3561 17980 3625 17984
rect 3561 17924 3565 17980
rect 3565 17924 3621 17980
rect 3621 17924 3625 17980
rect 3561 17920 3625 17924
rect 3641 17980 3705 17984
rect 3641 17924 3645 17980
rect 3645 17924 3701 17980
rect 3701 17924 3705 17980
rect 3641 17920 3705 17924
rect 8300 17980 8364 17984
rect 8300 17924 8304 17980
rect 8304 17924 8360 17980
rect 8360 17924 8364 17980
rect 8300 17920 8364 17924
rect 8380 17980 8444 17984
rect 8380 17924 8384 17980
rect 8384 17924 8440 17980
rect 8440 17924 8444 17980
rect 8380 17920 8444 17924
rect 8460 17980 8524 17984
rect 8460 17924 8464 17980
rect 8464 17924 8520 17980
rect 8520 17924 8524 17980
rect 8460 17920 8524 17924
rect 8540 17980 8604 17984
rect 8540 17924 8544 17980
rect 8544 17924 8600 17980
rect 8600 17924 8604 17980
rect 8540 17920 8604 17924
rect 13199 17980 13263 17984
rect 13199 17924 13203 17980
rect 13203 17924 13259 17980
rect 13259 17924 13263 17980
rect 13199 17920 13263 17924
rect 13279 17980 13343 17984
rect 13279 17924 13283 17980
rect 13283 17924 13339 17980
rect 13339 17924 13343 17980
rect 13279 17920 13343 17924
rect 13359 17980 13423 17984
rect 13359 17924 13363 17980
rect 13363 17924 13419 17980
rect 13419 17924 13423 17980
rect 13359 17920 13423 17924
rect 13439 17980 13503 17984
rect 13439 17924 13443 17980
rect 13443 17924 13499 17980
rect 13499 17924 13503 17980
rect 13439 17920 13503 17924
rect 18098 17980 18162 17984
rect 18098 17924 18102 17980
rect 18102 17924 18158 17980
rect 18158 17924 18162 17980
rect 18098 17920 18162 17924
rect 18178 17980 18242 17984
rect 18178 17924 18182 17980
rect 18182 17924 18238 17980
rect 18238 17924 18242 17980
rect 18178 17920 18242 17924
rect 18258 17980 18322 17984
rect 18258 17924 18262 17980
rect 18262 17924 18318 17980
rect 18318 17924 18322 17980
rect 18258 17920 18322 17924
rect 18338 17980 18402 17984
rect 18338 17924 18342 17980
rect 18342 17924 18398 17980
rect 18398 17924 18402 17980
rect 18338 17920 18402 17924
rect 5850 17436 5914 17440
rect 5850 17380 5854 17436
rect 5854 17380 5910 17436
rect 5910 17380 5914 17436
rect 5850 17376 5914 17380
rect 5930 17436 5994 17440
rect 5930 17380 5934 17436
rect 5934 17380 5990 17436
rect 5990 17380 5994 17436
rect 5930 17376 5994 17380
rect 6010 17436 6074 17440
rect 6010 17380 6014 17436
rect 6014 17380 6070 17436
rect 6070 17380 6074 17436
rect 6010 17376 6074 17380
rect 6090 17436 6154 17440
rect 6090 17380 6094 17436
rect 6094 17380 6150 17436
rect 6150 17380 6154 17436
rect 6090 17376 6154 17380
rect 10749 17436 10813 17440
rect 10749 17380 10753 17436
rect 10753 17380 10809 17436
rect 10809 17380 10813 17436
rect 10749 17376 10813 17380
rect 10829 17436 10893 17440
rect 10829 17380 10833 17436
rect 10833 17380 10889 17436
rect 10889 17380 10893 17436
rect 10829 17376 10893 17380
rect 10909 17436 10973 17440
rect 10909 17380 10913 17436
rect 10913 17380 10969 17436
rect 10969 17380 10973 17436
rect 10909 17376 10973 17380
rect 10989 17436 11053 17440
rect 10989 17380 10993 17436
rect 10993 17380 11049 17436
rect 11049 17380 11053 17436
rect 10989 17376 11053 17380
rect 15648 17436 15712 17440
rect 15648 17380 15652 17436
rect 15652 17380 15708 17436
rect 15708 17380 15712 17436
rect 15648 17376 15712 17380
rect 15728 17436 15792 17440
rect 15728 17380 15732 17436
rect 15732 17380 15788 17436
rect 15788 17380 15792 17436
rect 15728 17376 15792 17380
rect 15808 17436 15872 17440
rect 15808 17380 15812 17436
rect 15812 17380 15868 17436
rect 15868 17380 15872 17436
rect 15808 17376 15872 17380
rect 15888 17436 15952 17440
rect 15888 17380 15892 17436
rect 15892 17380 15948 17436
rect 15948 17380 15952 17436
rect 15888 17376 15952 17380
rect 20547 17436 20611 17440
rect 20547 17380 20551 17436
rect 20551 17380 20607 17436
rect 20607 17380 20611 17436
rect 20547 17376 20611 17380
rect 20627 17436 20691 17440
rect 20627 17380 20631 17436
rect 20631 17380 20687 17436
rect 20687 17380 20691 17436
rect 20627 17376 20691 17380
rect 20707 17436 20771 17440
rect 20707 17380 20711 17436
rect 20711 17380 20767 17436
rect 20767 17380 20771 17436
rect 20707 17376 20771 17380
rect 20787 17436 20851 17440
rect 20787 17380 20791 17436
rect 20791 17380 20847 17436
rect 20847 17380 20851 17436
rect 20787 17376 20851 17380
rect 3401 16892 3465 16896
rect 3401 16836 3405 16892
rect 3405 16836 3461 16892
rect 3461 16836 3465 16892
rect 3401 16832 3465 16836
rect 3481 16892 3545 16896
rect 3481 16836 3485 16892
rect 3485 16836 3541 16892
rect 3541 16836 3545 16892
rect 3481 16832 3545 16836
rect 3561 16892 3625 16896
rect 3561 16836 3565 16892
rect 3565 16836 3621 16892
rect 3621 16836 3625 16892
rect 3561 16832 3625 16836
rect 3641 16892 3705 16896
rect 3641 16836 3645 16892
rect 3645 16836 3701 16892
rect 3701 16836 3705 16892
rect 3641 16832 3705 16836
rect 8300 16892 8364 16896
rect 8300 16836 8304 16892
rect 8304 16836 8360 16892
rect 8360 16836 8364 16892
rect 8300 16832 8364 16836
rect 8380 16892 8444 16896
rect 8380 16836 8384 16892
rect 8384 16836 8440 16892
rect 8440 16836 8444 16892
rect 8380 16832 8444 16836
rect 8460 16892 8524 16896
rect 8460 16836 8464 16892
rect 8464 16836 8520 16892
rect 8520 16836 8524 16892
rect 8460 16832 8524 16836
rect 8540 16892 8604 16896
rect 8540 16836 8544 16892
rect 8544 16836 8600 16892
rect 8600 16836 8604 16892
rect 8540 16832 8604 16836
rect 13199 16892 13263 16896
rect 13199 16836 13203 16892
rect 13203 16836 13259 16892
rect 13259 16836 13263 16892
rect 13199 16832 13263 16836
rect 13279 16892 13343 16896
rect 13279 16836 13283 16892
rect 13283 16836 13339 16892
rect 13339 16836 13343 16892
rect 13279 16832 13343 16836
rect 13359 16892 13423 16896
rect 13359 16836 13363 16892
rect 13363 16836 13419 16892
rect 13419 16836 13423 16892
rect 13359 16832 13423 16836
rect 13439 16892 13503 16896
rect 13439 16836 13443 16892
rect 13443 16836 13499 16892
rect 13499 16836 13503 16892
rect 13439 16832 13503 16836
rect 18098 16892 18162 16896
rect 18098 16836 18102 16892
rect 18102 16836 18158 16892
rect 18158 16836 18162 16892
rect 18098 16832 18162 16836
rect 18178 16892 18242 16896
rect 18178 16836 18182 16892
rect 18182 16836 18238 16892
rect 18238 16836 18242 16892
rect 18178 16832 18242 16836
rect 18258 16892 18322 16896
rect 18258 16836 18262 16892
rect 18262 16836 18318 16892
rect 18318 16836 18322 16892
rect 18258 16832 18322 16836
rect 18338 16892 18402 16896
rect 18338 16836 18342 16892
rect 18342 16836 18398 16892
rect 18398 16836 18402 16892
rect 18338 16832 18402 16836
rect 5850 16348 5914 16352
rect 5850 16292 5854 16348
rect 5854 16292 5910 16348
rect 5910 16292 5914 16348
rect 5850 16288 5914 16292
rect 5930 16348 5994 16352
rect 5930 16292 5934 16348
rect 5934 16292 5990 16348
rect 5990 16292 5994 16348
rect 5930 16288 5994 16292
rect 6010 16348 6074 16352
rect 6010 16292 6014 16348
rect 6014 16292 6070 16348
rect 6070 16292 6074 16348
rect 6010 16288 6074 16292
rect 6090 16348 6154 16352
rect 6090 16292 6094 16348
rect 6094 16292 6150 16348
rect 6150 16292 6154 16348
rect 6090 16288 6154 16292
rect 10749 16348 10813 16352
rect 10749 16292 10753 16348
rect 10753 16292 10809 16348
rect 10809 16292 10813 16348
rect 10749 16288 10813 16292
rect 10829 16348 10893 16352
rect 10829 16292 10833 16348
rect 10833 16292 10889 16348
rect 10889 16292 10893 16348
rect 10829 16288 10893 16292
rect 10909 16348 10973 16352
rect 10909 16292 10913 16348
rect 10913 16292 10969 16348
rect 10969 16292 10973 16348
rect 10909 16288 10973 16292
rect 10989 16348 11053 16352
rect 10989 16292 10993 16348
rect 10993 16292 11049 16348
rect 11049 16292 11053 16348
rect 10989 16288 11053 16292
rect 15648 16348 15712 16352
rect 15648 16292 15652 16348
rect 15652 16292 15708 16348
rect 15708 16292 15712 16348
rect 15648 16288 15712 16292
rect 15728 16348 15792 16352
rect 15728 16292 15732 16348
rect 15732 16292 15788 16348
rect 15788 16292 15792 16348
rect 15728 16288 15792 16292
rect 15808 16348 15872 16352
rect 15808 16292 15812 16348
rect 15812 16292 15868 16348
rect 15868 16292 15872 16348
rect 15808 16288 15872 16292
rect 15888 16348 15952 16352
rect 15888 16292 15892 16348
rect 15892 16292 15948 16348
rect 15948 16292 15952 16348
rect 15888 16288 15952 16292
rect 20547 16348 20611 16352
rect 20547 16292 20551 16348
rect 20551 16292 20607 16348
rect 20607 16292 20611 16348
rect 20547 16288 20611 16292
rect 20627 16348 20691 16352
rect 20627 16292 20631 16348
rect 20631 16292 20687 16348
rect 20687 16292 20691 16348
rect 20627 16288 20691 16292
rect 20707 16348 20771 16352
rect 20707 16292 20711 16348
rect 20711 16292 20767 16348
rect 20767 16292 20771 16348
rect 20707 16288 20771 16292
rect 20787 16348 20851 16352
rect 20787 16292 20791 16348
rect 20791 16292 20847 16348
rect 20847 16292 20851 16348
rect 20787 16288 20851 16292
rect 3401 15804 3465 15808
rect 3401 15748 3405 15804
rect 3405 15748 3461 15804
rect 3461 15748 3465 15804
rect 3401 15744 3465 15748
rect 3481 15804 3545 15808
rect 3481 15748 3485 15804
rect 3485 15748 3541 15804
rect 3541 15748 3545 15804
rect 3481 15744 3545 15748
rect 3561 15804 3625 15808
rect 3561 15748 3565 15804
rect 3565 15748 3621 15804
rect 3621 15748 3625 15804
rect 3561 15744 3625 15748
rect 3641 15804 3705 15808
rect 3641 15748 3645 15804
rect 3645 15748 3701 15804
rect 3701 15748 3705 15804
rect 3641 15744 3705 15748
rect 8300 15804 8364 15808
rect 8300 15748 8304 15804
rect 8304 15748 8360 15804
rect 8360 15748 8364 15804
rect 8300 15744 8364 15748
rect 8380 15804 8444 15808
rect 8380 15748 8384 15804
rect 8384 15748 8440 15804
rect 8440 15748 8444 15804
rect 8380 15744 8444 15748
rect 8460 15804 8524 15808
rect 8460 15748 8464 15804
rect 8464 15748 8520 15804
rect 8520 15748 8524 15804
rect 8460 15744 8524 15748
rect 8540 15804 8604 15808
rect 8540 15748 8544 15804
rect 8544 15748 8600 15804
rect 8600 15748 8604 15804
rect 8540 15744 8604 15748
rect 13199 15804 13263 15808
rect 13199 15748 13203 15804
rect 13203 15748 13259 15804
rect 13259 15748 13263 15804
rect 13199 15744 13263 15748
rect 13279 15804 13343 15808
rect 13279 15748 13283 15804
rect 13283 15748 13339 15804
rect 13339 15748 13343 15804
rect 13279 15744 13343 15748
rect 13359 15804 13423 15808
rect 13359 15748 13363 15804
rect 13363 15748 13419 15804
rect 13419 15748 13423 15804
rect 13359 15744 13423 15748
rect 13439 15804 13503 15808
rect 13439 15748 13443 15804
rect 13443 15748 13499 15804
rect 13499 15748 13503 15804
rect 13439 15744 13503 15748
rect 18098 15804 18162 15808
rect 18098 15748 18102 15804
rect 18102 15748 18158 15804
rect 18158 15748 18162 15804
rect 18098 15744 18162 15748
rect 18178 15804 18242 15808
rect 18178 15748 18182 15804
rect 18182 15748 18238 15804
rect 18238 15748 18242 15804
rect 18178 15744 18242 15748
rect 18258 15804 18322 15808
rect 18258 15748 18262 15804
rect 18262 15748 18318 15804
rect 18318 15748 18322 15804
rect 18258 15744 18322 15748
rect 18338 15804 18402 15808
rect 18338 15748 18342 15804
rect 18342 15748 18398 15804
rect 18398 15748 18402 15804
rect 18338 15744 18402 15748
rect 5850 15260 5914 15264
rect 5850 15204 5854 15260
rect 5854 15204 5910 15260
rect 5910 15204 5914 15260
rect 5850 15200 5914 15204
rect 5930 15260 5994 15264
rect 5930 15204 5934 15260
rect 5934 15204 5990 15260
rect 5990 15204 5994 15260
rect 5930 15200 5994 15204
rect 6010 15260 6074 15264
rect 6010 15204 6014 15260
rect 6014 15204 6070 15260
rect 6070 15204 6074 15260
rect 6010 15200 6074 15204
rect 6090 15260 6154 15264
rect 6090 15204 6094 15260
rect 6094 15204 6150 15260
rect 6150 15204 6154 15260
rect 6090 15200 6154 15204
rect 10749 15260 10813 15264
rect 10749 15204 10753 15260
rect 10753 15204 10809 15260
rect 10809 15204 10813 15260
rect 10749 15200 10813 15204
rect 10829 15260 10893 15264
rect 10829 15204 10833 15260
rect 10833 15204 10889 15260
rect 10889 15204 10893 15260
rect 10829 15200 10893 15204
rect 10909 15260 10973 15264
rect 10909 15204 10913 15260
rect 10913 15204 10969 15260
rect 10969 15204 10973 15260
rect 10909 15200 10973 15204
rect 10989 15260 11053 15264
rect 10989 15204 10993 15260
rect 10993 15204 11049 15260
rect 11049 15204 11053 15260
rect 10989 15200 11053 15204
rect 15648 15260 15712 15264
rect 15648 15204 15652 15260
rect 15652 15204 15708 15260
rect 15708 15204 15712 15260
rect 15648 15200 15712 15204
rect 15728 15260 15792 15264
rect 15728 15204 15732 15260
rect 15732 15204 15788 15260
rect 15788 15204 15792 15260
rect 15728 15200 15792 15204
rect 15808 15260 15872 15264
rect 15808 15204 15812 15260
rect 15812 15204 15868 15260
rect 15868 15204 15872 15260
rect 15808 15200 15872 15204
rect 15888 15260 15952 15264
rect 15888 15204 15892 15260
rect 15892 15204 15948 15260
rect 15948 15204 15952 15260
rect 15888 15200 15952 15204
rect 20547 15260 20611 15264
rect 20547 15204 20551 15260
rect 20551 15204 20607 15260
rect 20607 15204 20611 15260
rect 20547 15200 20611 15204
rect 20627 15260 20691 15264
rect 20627 15204 20631 15260
rect 20631 15204 20687 15260
rect 20687 15204 20691 15260
rect 20627 15200 20691 15204
rect 20707 15260 20771 15264
rect 20707 15204 20711 15260
rect 20711 15204 20767 15260
rect 20767 15204 20771 15260
rect 20707 15200 20771 15204
rect 20787 15260 20851 15264
rect 20787 15204 20791 15260
rect 20791 15204 20847 15260
rect 20847 15204 20851 15260
rect 20787 15200 20851 15204
rect 3401 14716 3465 14720
rect 3401 14660 3405 14716
rect 3405 14660 3461 14716
rect 3461 14660 3465 14716
rect 3401 14656 3465 14660
rect 3481 14716 3545 14720
rect 3481 14660 3485 14716
rect 3485 14660 3541 14716
rect 3541 14660 3545 14716
rect 3481 14656 3545 14660
rect 3561 14716 3625 14720
rect 3561 14660 3565 14716
rect 3565 14660 3621 14716
rect 3621 14660 3625 14716
rect 3561 14656 3625 14660
rect 3641 14716 3705 14720
rect 3641 14660 3645 14716
rect 3645 14660 3701 14716
rect 3701 14660 3705 14716
rect 3641 14656 3705 14660
rect 8300 14716 8364 14720
rect 8300 14660 8304 14716
rect 8304 14660 8360 14716
rect 8360 14660 8364 14716
rect 8300 14656 8364 14660
rect 8380 14716 8444 14720
rect 8380 14660 8384 14716
rect 8384 14660 8440 14716
rect 8440 14660 8444 14716
rect 8380 14656 8444 14660
rect 8460 14716 8524 14720
rect 8460 14660 8464 14716
rect 8464 14660 8520 14716
rect 8520 14660 8524 14716
rect 8460 14656 8524 14660
rect 8540 14716 8604 14720
rect 8540 14660 8544 14716
rect 8544 14660 8600 14716
rect 8600 14660 8604 14716
rect 8540 14656 8604 14660
rect 13199 14716 13263 14720
rect 13199 14660 13203 14716
rect 13203 14660 13259 14716
rect 13259 14660 13263 14716
rect 13199 14656 13263 14660
rect 13279 14716 13343 14720
rect 13279 14660 13283 14716
rect 13283 14660 13339 14716
rect 13339 14660 13343 14716
rect 13279 14656 13343 14660
rect 13359 14716 13423 14720
rect 13359 14660 13363 14716
rect 13363 14660 13419 14716
rect 13419 14660 13423 14716
rect 13359 14656 13423 14660
rect 13439 14716 13503 14720
rect 13439 14660 13443 14716
rect 13443 14660 13499 14716
rect 13499 14660 13503 14716
rect 13439 14656 13503 14660
rect 18098 14716 18162 14720
rect 18098 14660 18102 14716
rect 18102 14660 18158 14716
rect 18158 14660 18162 14716
rect 18098 14656 18162 14660
rect 18178 14716 18242 14720
rect 18178 14660 18182 14716
rect 18182 14660 18238 14716
rect 18238 14660 18242 14716
rect 18178 14656 18242 14660
rect 18258 14716 18322 14720
rect 18258 14660 18262 14716
rect 18262 14660 18318 14716
rect 18318 14660 18322 14716
rect 18258 14656 18322 14660
rect 18338 14716 18402 14720
rect 18338 14660 18342 14716
rect 18342 14660 18398 14716
rect 18398 14660 18402 14716
rect 18338 14656 18402 14660
rect 5850 14172 5914 14176
rect 5850 14116 5854 14172
rect 5854 14116 5910 14172
rect 5910 14116 5914 14172
rect 5850 14112 5914 14116
rect 5930 14172 5994 14176
rect 5930 14116 5934 14172
rect 5934 14116 5990 14172
rect 5990 14116 5994 14172
rect 5930 14112 5994 14116
rect 6010 14172 6074 14176
rect 6010 14116 6014 14172
rect 6014 14116 6070 14172
rect 6070 14116 6074 14172
rect 6010 14112 6074 14116
rect 6090 14172 6154 14176
rect 6090 14116 6094 14172
rect 6094 14116 6150 14172
rect 6150 14116 6154 14172
rect 6090 14112 6154 14116
rect 10749 14172 10813 14176
rect 10749 14116 10753 14172
rect 10753 14116 10809 14172
rect 10809 14116 10813 14172
rect 10749 14112 10813 14116
rect 10829 14172 10893 14176
rect 10829 14116 10833 14172
rect 10833 14116 10889 14172
rect 10889 14116 10893 14172
rect 10829 14112 10893 14116
rect 10909 14172 10973 14176
rect 10909 14116 10913 14172
rect 10913 14116 10969 14172
rect 10969 14116 10973 14172
rect 10909 14112 10973 14116
rect 10989 14172 11053 14176
rect 10989 14116 10993 14172
rect 10993 14116 11049 14172
rect 11049 14116 11053 14172
rect 10989 14112 11053 14116
rect 15648 14172 15712 14176
rect 15648 14116 15652 14172
rect 15652 14116 15708 14172
rect 15708 14116 15712 14172
rect 15648 14112 15712 14116
rect 15728 14172 15792 14176
rect 15728 14116 15732 14172
rect 15732 14116 15788 14172
rect 15788 14116 15792 14172
rect 15728 14112 15792 14116
rect 15808 14172 15872 14176
rect 15808 14116 15812 14172
rect 15812 14116 15868 14172
rect 15868 14116 15872 14172
rect 15808 14112 15872 14116
rect 15888 14172 15952 14176
rect 15888 14116 15892 14172
rect 15892 14116 15948 14172
rect 15948 14116 15952 14172
rect 15888 14112 15952 14116
rect 20547 14172 20611 14176
rect 20547 14116 20551 14172
rect 20551 14116 20607 14172
rect 20607 14116 20611 14172
rect 20547 14112 20611 14116
rect 20627 14172 20691 14176
rect 20627 14116 20631 14172
rect 20631 14116 20687 14172
rect 20687 14116 20691 14172
rect 20627 14112 20691 14116
rect 20707 14172 20771 14176
rect 20707 14116 20711 14172
rect 20711 14116 20767 14172
rect 20767 14116 20771 14172
rect 20707 14112 20771 14116
rect 20787 14172 20851 14176
rect 20787 14116 20791 14172
rect 20791 14116 20847 14172
rect 20847 14116 20851 14172
rect 20787 14112 20851 14116
rect 3401 13628 3465 13632
rect 3401 13572 3405 13628
rect 3405 13572 3461 13628
rect 3461 13572 3465 13628
rect 3401 13568 3465 13572
rect 3481 13628 3545 13632
rect 3481 13572 3485 13628
rect 3485 13572 3541 13628
rect 3541 13572 3545 13628
rect 3481 13568 3545 13572
rect 3561 13628 3625 13632
rect 3561 13572 3565 13628
rect 3565 13572 3621 13628
rect 3621 13572 3625 13628
rect 3561 13568 3625 13572
rect 3641 13628 3705 13632
rect 3641 13572 3645 13628
rect 3645 13572 3701 13628
rect 3701 13572 3705 13628
rect 3641 13568 3705 13572
rect 8300 13628 8364 13632
rect 8300 13572 8304 13628
rect 8304 13572 8360 13628
rect 8360 13572 8364 13628
rect 8300 13568 8364 13572
rect 8380 13628 8444 13632
rect 8380 13572 8384 13628
rect 8384 13572 8440 13628
rect 8440 13572 8444 13628
rect 8380 13568 8444 13572
rect 8460 13628 8524 13632
rect 8460 13572 8464 13628
rect 8464 13572 8520 13628
rect 8520 13572 8524 13628
rect 8460 13568 8524 13572
rect 8540 13628 8604 13632
rect 8540 13572 8544 13628
rect 8544 13572 8600 13628
rect 8600 13572 8604 13628
rect 8540 13568 8604 13572
rect 13199 13628 13263 13632
rect 13199 13572 13203 13628
rect 13203 13572 13259 13628
rect 13259 13572 13263 13628
rect 13199 13568 13263 13572
rect 13279 13628 13343 13632
rect 13279 13572 13283 13628
rect 13283 13572 13339 13628
rect 13339 13572 13343 13628
rect 13279 13568 13343 13572
rect 13359 13628 13423 13632
rect 13359 13572 13363 13628
rect 13363 13572 13419 13628
rect 13419 13572 13423 13628
rect 13359 13568 13423 13572
rect 13439 13628 13503 13632
rect 13439 13572 13443 13628
rect 13443 13572 13499 13628
rect 13499 13572 13503 13628
rect 13439 13568 13503 13572
rect 18098 13628 18162 13632
rect 18098 13572 18102 13628
rect 18102 13572 18158 13628
rect 18158 13572 18162 13628
rect 18098 13568 18162 13572
rect 18178 13628 18242 13632
rect 18178 13572 18182 13628
rect 18182 13572 18238 13628
rect 18238 13572 18242 13628
rect 18178 13568 18242 13572
rect 18258 13628 18322 13632
rect 18258 13572 18262 13628
rect 18262 13572 18318 13628
rect 18318 13572 18322 13628
rect 18258 13568 18322 13572
rect 18338 13628 18402 13632
rect 18338 13572 18342 13628
rect 18342 13572 18398 13628
rect 18398 13572 18402 13628
rect 18338 13568 18402 13572
rect 5850 13084 5914 13088
rect 5850 13028 5854 13084
rect 5854 13028 5910 13084
rect 5910 13028 5914 13084
rect 5850 13024 5914 13028
rect 5930 13084 5994 13088
rect 5930 13028 5934 13084
rect 5934 13028 5990 13084
rect 5990 13028 5994 13084
rect 5930 13024 5994 13028
rect 6010 13084 6074 13088
rect 6010 13028 6014 13084
rect 6014 13028 6070 13084
rect 6070 13028 6074 13084
rect 6010 13024 6074 13028
rect 6090 13084 6154 13088
rect 6090 13028 6094 13084
rect 6094 13028 6150 13084
rect 6150 13028 6154 13084
rect 6090 13024 6154 13028
rect 10749 13084 10813 13088
rect 10749 13028 10753 13084
rect 10753 13028 10809 13084
rect 10809 13028 10813 13084
rect 10749 13024 10813 13028
rect 10829 13084 10893 13088
rect 10829 13028 10833 13084
rect 10833 13028 10889 13084
rect 10889 13028 10893 13084
rect 10829 13024 10893 13028
rect 10909 13084 10973 13088
rect 10909 13028 10913 13084
rect 10913 13028 10969 13084
rect 10969 13028 10973 13084
rect 10909 13024 10973 13028
rect 10989 13084 11053 13088
rect 10989 13028 10993 13084
rect 10993 13028 11049 13084
rect 11049 13028 11053 13084
rect 10989 13024 11053 13028
rect 15648 13084 15712 13088
rect 15648 13028 15652 13084
rect 15652 13028 15708 13084
rect 15708 13028 15712 13084
rect 15648 13024 15712 13028
rect 15728 13084 15792 13088
rect 15728 13028 15732 13084
rect 15732 13028 15788 13084
rect 15788 13028 15792 13084
rect 15728 13024 15792 13028
rect 15808 13084 15872 13088
rect 15808 13028 15812 13084
rect 15812 13028 15868 13084
rect 15868 13028 15872 13084
rect 15808 13024 15872 13028
rect 15888 13084 15952 13088
rect 15888 13028 15892 13084
rect 15892 13028 15948 13084
rect 15948 13028 15952 13084
rect 15888 13024 15952 13028
rect 20547 13084 20611 13088
rect 20547 13028 20551 13084
rect 20551 13028 20607 13084
rect 20607 13028 20611 13084
rect 20547 13024 20611 13028
rect 20627 13084 20691 13088
rect 20627 13028 20631 13084
rect 20631 13028 20687 13084
rect 20687 13028 20691 13084
rect 20627 13024 20691 13028
rect 20707 13084 20771 13088
rect 20707 13028 20711 13084
rect 20711 13028 20767 13084
rect 20767 13028 20771 13084
rect 20707 13024 20771 13028
rect 20787 13084 20851 13088
rect 20787 13028 20791 13084
rect 20791 13028 20847 13084
rect 20847 13028 20851 13084
rect 20787 13024 20851 13028
rect 3401 12540 3465 12544
rect 3401 12484 3405 12540
rect 3405 12484 3461 12540
rect 3461 12484 3465 12540
rect 3401 12480 3465 12484
rect 3481 12540 3545 12544
rect 3481 12484 3485 12540
rect 3485 12484 3541 12540
rect 3541 12484 3545 12540
rect 3481 12480 3545 12484
rect 3561 12540 3625 12544
rect 3561 12484 3565 12540
rect 3565 12484 3621 12540
rect 3621 12484 3625 12540
rect 3561 12480 3625 12484
rect 3641 12540 3705 12544
rect 3641 12484 3645 12540
rect 3645 12484 3701 12540
rect 3701 12484 3705 12540
rect 3641 12480 3705 12484
rect 8300 12540 8364 12544
rect 8300 12484 8304 12540
rect 8304 12484 8360 12540
rect 8360 12484 8364 12540
rect 8300 12480 8364 12484
rect 8380 12540 8444 12544
rect 8380 12484 8384 12540
rect 8384 12484 8440 12540
rect 8440 12484 8444 12540
rect 8380 12480 8444 12484
rect 8460 12540 8524 12544
rect 8460 12484 8464 12540
rect 8464 12484 8520 12540
rect 8520 12484 8524 12540
rect 8460 12480 8524 12484
rect 8540 12540 8604 12544
rect 8540 12484 8544 12540
rect 8544 12484 8600 12540
rect 8600 12484 8604 12540
rect 8540 12480 8604 12484
rect 13199 12540 13263 12544
rect 13199 12484 13203 12540
rect 13203 12484 13259 12540
rect 13259 12484 13263 12540
rect 13199 12480 13263 12484
rect 13279 12540 13343 12544
rect 13279 12484 13283 12540
rect 13283 12484 13339 12540
rect 13339 12484 13343 12540
rect 13279 12480 13343 12484
rect 13359 12540 13423 12544
rect 13359 12484 13363 12540
rect 13363 12484 13419 12540
rect 13419 12484 13423 12540
rect 13359 12480 13423 12484
rect 13439 12540 13503 12544
rect 13439 12484 13443 12540
rect 13443 12484 13499 12540
rect 13499 12484 13503 12540
rect 13439 12480 13503 12484
rect 18098 12540 18162 12544
rect 18098 12484 18102 12540
rect 18102 12484 18158 12540
rect 18158 12484 18162 12540
rect 18098 12480 18162 12484
rect 18178 12540 18242 12544
rect 18178 12484 18182 12540
rect 18182 12484 18238 12540
rect 18238 12484 18242 12540
rect 18178 12480 18242 12484
rect 18258 12540 18322 12544
rect 18258 12484 18262 12540
rect 18262 12484 18318 12540
rect 18318 12484 18322 12540
rect 18258 12480 18322 12484
rect 18338 12540 18402 12544
rect 18338 12484 18342 12540
rect 18342 12484 18398 12540
rect 18398 12484 18402 12540
rect 18338 12480 18402 12484
rect 5850 11996 5914 12000
rect 5850 11940 5854 11996
rect 5854 11940 5910 11996
rect 5910 11940 5914 11996
rect 5850 11936 5914 11940
rect 5930 11996 5994 12000
rect 5930 11940 5934 11996
rect 5934 11940 5990 11996
rect 5990 11940 5994 11996
rect 5930 11936 5994 11940
rect 6010 11996 6074 12000
rect 6010 11940 6014 11996
rect 6014 11940 6070 11996
rect 6070 11940 6074 11996
rect 6010 11936 6074 11940
rect 6090 11996 6154 12000
rect 6090 11940 6094 11996
rect 6094 11940 6150 11996
rect 6150 11940 6154 11996
rect 6090 11936 6154 11940
rect 10749 11996 10813 12000
rect 10749 11940 10753 11996
rect 10753 11940 10809 11996
rect 10809 11940 10813 11996
rect 10749 11936 10813 11940
rect 10829 11996 10893 12000
rect 10829 11940 10833 11996
rect 10833 11940 10889 11996
rect 10889 11940 10893 11996
rect 10829 11936 10893 11940
rect 10909 11996 10973 12000
rect 10909 11940 10913 11996
rect 10913 11940 10969 11996
rect 10969 11940 10973 11996
rect 10909 11936 10973 11940
rect 10989 11996 11053 12000
rect 10989 11940 10993 11996
rect 10993 11940 11049 11996
rect 11049 11940 11053 11996
rect 10989 11936 11053 11940
rect 15648 11996 15712 12000
rect 15648 11940 15652 11996
rect 15652 11940 15708 11996
rect 15708 11940 15712 11996
rect 15648 11936 15712 11940
rect 15728 11996 15792 12000
rect 15728 11940 15732 11996
rect 15732 11940 15788 11996
rect 15788 11940 15792 11996
rect 15728 11936 15792 11940
rect 15808 11996 15872 12000
rect 15808 11940 15812 11996
rect 15812 11940 15868 11996
rect 15868 11940 15872 11996
rect 15808 11936 15872 11940
rect 15888 11996 15952 12000
rect 15888 11940 15892 11996
rect 15892 11940 15948 11996
rect 15948 11940 15952 11996
rect 15888 11936 15952 11940
rect 20547 11996 20611 12000
rect 20547 11940 20551 11996
rect 20551 11940 20607 11996
rect 20607 11940 20611 11996
rect 20547 11936 20611 11940
rect 20627 11996 20691 12000
rect 20627 11940 20631 11996
rect 20631 11940 20687 11996
rect 20687 11940 20691 11996
rect 20627 11936 20691 11940
rect 20707 11996 20771 12000
rect 20707 11940 20711 11996
rect 20711 11940 20767 11996
rect 20767 11940 20771 11996
rect 20707 11936 20771 11940
rect 20787 11996 20851 12000
rect 20787 11940 20791 11996
rect 20791 11940 20847 11996
rect 20847 11940 20851 11996
rect 20787 11936 20851 11940
rect 3401 11452 3465 11456
rect 3401 11396 3405 11452
rect 3405 11396 3461 11452
rect 3461 11396 3465 11452
rect 3401 11392 3465 11396
rect 3481 11452 3545 11456
rect 3481 11396 3485 11452
rect 3485 11396 3541 11452
rect 3541 11396 3545 11452
rect 3481 11392 3545 11396
rect 3561 11452 3625 11456
rect 3561 11396 3565 11452
rect 3565 11396 3621 11452
rect 3621 11396 3625 11452
rect 3561 11392 3625 11396
rect 3641 11452 3705 11456
rect 3641 11396 3645 11452
rect 3645 11396 3701 11452
rect 3701 11396 3705 11452
rect 3641 11392 3705 11396
rect 8300 11452 8364 11456
rect 8300 11396 8304 11452
rect 8304 11396 8360 11452
rect 8360 11396 8364 11452
rect 8300 11392 8364 11396
rect 8380 11452 8444 11456
rect 8380 11396 8384 11452
rect 8384 11396 8440 11452
rect 8440 11396 8444 11452
rect 8380 11392 8444 11396
rect 8460 11452 8524 11456
rect 8460 11396 8464 11452
rect 8464 11396 8520 11452
rect 8520 11396 8524 11452
rect 8460 11392 8524 11396
rect 8540 11452 8604 11456
rect 8540 11396 8544 11452
rect 8544 11396 8600 11452
rect 8600 11396 8604 11452
rect 8540 11392 8604 11396
rect 13199 11452 13263 11456
rect 13199 11396 13203 11452
rect 13203 11396 13259 11452
rect 13259 11396 13263 11452
rect 13199 11392 13263 11396
rect 13279 11452 13343 11456
rect 13279 11396 13283 11452
rect 13283 11396 13339 11452
rect 13339 11396 13343 11452
rect 13279 11392 13343 11396
rect 13359 11452 13423 11456
rect 13359 11396 13363 11452
rect 13363 11396 13419 11452
rect 13419 11396 13423 11452
rect 13359 11392 13423 11396
rect 13439 11452 13503 11456
rect 13439 11396 13443 11452
rect 13443 11396 13499 11452
rect 13499 11396 13503 11452
rect 13439 11392 13503 11396
rect 18098 11452 18162 11456
rect 18098 11396 18102 11452
rect 18102 11396 18158 11452
rect 18158 11396 18162 11452
rect 18098 11392 18162 11396
rect 18178 11452 18242 11456
rect 18178 11396 18182 11452
rect 18182 11396 18238 11452
rect 18238 11396 18242 11452
rect 18178 11392 18242 11396
rect 18258 11452 18322 11456
rect 18258 11396 18262 11452
rect 18262 11396 18318 11452
rect 18318 11396 18322 11452
rect 18258 11392 18322 11396
rect 18338 11452 18402 11456
rect 18338 11396 18342 11452
rect 18342 11396 18398 11452
rect 18398 11396 18402 11452
rect 18338 11392 18402 11396
rect 5850 10908 5914 10912
rect 5850 10852 5854 10908
rect 5854 10852 5910 10908
rect 5910 10852 5914 10908
rect 5850 10848 5914 10852
rect 5930 10908 5994 10912
rect 5930 10852 5934 10908
rect 5934 10852 5990 10908
rect 5990 10852 5994 10908
rect 5930 10848 5994 10852
rect 6010 10908 6074 10912
rect 6010 10852 6014 10908
rect 6014 10852 6070 10908
rect 6070 10852 6074 10908
rect 6010 10848 6074 10852
rect 6090 10908 6154 10912
rect 6090 10852 6094 10908
rect 6094 10852 6150 10908
rect 6150 10852 6154 10908
rect 6090 10848 6154 10852
rect 10749 10908 10813 10912
rect 10749 10852 10753 10908
rect 10753 10852 10809 10908
rect 10809 10852 10813 10908
rect 10749 10848 10813 10852
rect 10829 10908 10893 10912
rect 10829 10852 10833 10908
rect 10833 10852 10889 10908
rect 10889 10852 10893 10908
rect 10829 10848 10893 10852
rect 10909 10908 10973 10912
rect 10909 10852 10913 10908
rect 10913 10852 10969 10908
rect 10969 10852 10973 10908
rect 10909 10848 10973 10852
rect 10989 10908 11053 10912
rect 10989 10852 10993 10908
rect 10993 10852 11049 10908
rect 11049 10852 11053 10908
rect 10989 10848 11053 10852
rect 15648 10908 15712 10912
rect 15648 10852 15652 10908
rect 15652 10852 15708 10908
rect 15708 10852 15712 10908
rect 15648 10848 15712 10852
rect 15728 10908 15792 10912
rect 15728 10852 15732 10908
rect 15732 10852 15788 10908
rect 15788 10852 15792 10908
rect 15728 10848 15792 10852
rect 15808 10908 15872 10912
rect 15808 10852 15812 10908
rect 15812 10852 15868 10908
rect 15868 10852 15872 10908
rect 15808 10848 15872 10852
rect 15888 10908 15952 10912
rect 15888 10852 15892 10908
rect 15892 10852 15948 10908
rect 15948 10852 15952 10908
rect 15888 10848 15952 10852
rect 20547 10908 20611 10912
rect 20547 10852 20551 10908
rect 20551 10852 20607 10908
rect 20607 10852 20611 10908
rect 20547 10848 20611 10852
rect 20627 10908 20691 10912
rect 20627 10852 20631 10908
rect 20631 10852 20687 10908
rect 20687 10852 20691 10908
rect 20627 10848 20691 10852
rect 20707 10908 20771 10912
rect 20707 10852 20711 10908
rect 20711 10852 20767 10908
rect 20767 10852 20771 10908
rect 20707 10848 20771 10852
rect 20787 10908 20851 10912
rect 20787 10852 20791 10908
rect 20791 10852 20847 10908
rect 20847 10852 20851 10908
rect 20787 10848 20851 10852
rect 3401 10364 3465 10368
rect 3401 10308 3405 10364
rect 3405 10308 3461 10364
rect 3461 10308 3465 10364
rect 3401 10304 3465 10308
rect 3481 10364 3545 10368
rect 3481 10308 3485 10364
rect 3485 10308 3541 10364
rect 3541 10308 3545 10364
rect 3481 10304 3545 10308
rect 3561 10364 3625 10368
rect 3561 10308 3565 10364
rect 3565 10308 3621 10364
rect 3621 10308 3625 10364
rect 3561 10304 3625 10308
rect 3641 10364 3705 10368
rect 3641 10308 3645 10364
rect 3645 10308 3701 10364
rect 3701 10308 3705 10364
rect 3641 10304 3705 10308
rect 8300 10364 8364 10368
rect 8300 10308 8304 10364
rect 8304 10308 8360 10364
rect 8360 10308 8364 10364
rect 8300 10304 8364 10308
rect 8380 10364 8444 10368
rect 8380 10308 8384 10364
rect 8384 10308 8440 10364
rect 8440 10308 8444 10364
rect 8380 10304 8444 10308
rect 8460 10364 8524 10368
rect 8460 10308 8464 10364
rect 8464 10308 8520 10364
rect 8520 10308 8524 10364
rect 8460 10304 8524 10308
rect 8540 10364 8604 10368
rect 8540 10308 8544 10364
rect 8544 10308 8600 10364
rect 8600 10308 8604 10364
rect 8540 10304 8604 10308
rect 13199 10364 13263 10368
rect 13199 10308 13203 10364
rect 13203 10308 13259 10364
rect 13259 10308 13263 10364
rect 13199 10304 13263 10308
rect 13279 10364 13343 10368
rect 13279 10308 13283 10364
rect 13283 10308 13339 10364
rect 13339 10308 13343 10364
rect 13279 10304 13343 10308
rect 13359 10364 13423 10368
rect 13359 10308 13363 10364
rect 13363 10308 13419 10364
rect 13419 10308 13423 10364
rect 13359 10304 13423 10308
rect 13439 10364 13503 10368
rect 13439 10308 13443 10364
rect 13443 10308 13499 10364
rect 13499 10308 13503 10364
rect 13439 10304 13503 10308
rect 18098 10364 18162 10368
rect 18098 10308 18102 10364
rect 18102 10308 18158 10364
rect 18158 10308 18162 10364
rect 18098 10304 18162 10308
rect 18178 10364 18242 10368
rect 18178 10308 18182 10364
rect 18182 10308 18238 10364
rect 18238 10308 18242 10364
rect 18178 10304 18242 10308
rect 18258 10364 18322 10368
rect 18258 10308 18262 10364
rect 18262 10308 18318 10364
rect 18318 10308 18322 10364
rect 18258 10304 18322 10308
rect 18338 10364 18402 10368
rect 18338 10308 18342 10364
rect 18342 10308 18398 10364
rect 18398 10308 18402 10364
rect 18338 10304 18402 10308
rect 5850 9820 5914 9824
rect 5850 9764 5854 9820
rect 5854 9764 5910 9820
rect 5910 9764 5914 9820
rect 5850 9760 5914 9764
rect 5930 9820 5994 9824
rect 5930 9764 5934 9820
rect 5934 9764 5990 9820
rect 5990 9764 5994 9820
rect 5930 9760 5994 9764
rect 6010 9820 6074 9824
rect 6010 9764 6014 9820
rect 6014 9764 6070 9820
rect 6070 9764 6074 9820
rect 6010 9760 6074 9764
rect 6090 9820 6154 9824
rect 6090 9764 6094 9820
rect 6094 9764 6150 9820
rect 6150 9764 6154 9820
rect 6090 9760 6154 9764
rect 10749 9820 10813 9824
rect 10749 9764 10753 9820
rect 10753 9764 10809 9820
rect 10809 9764 10813 9820
rect 10749 9760 10813 9764
rect 10829 9820 10893 9824
rect 10829 9764 10833 9820
rect 10833 9764 10889 9820
rect 10889 9764 10893 9820
rect 10829 9760 10893 9764
rect 10909 9820 10973 9824
rect 10909 9764 10913 9820
rect 10913 9764 10969 9820
rect 10969 9764 10973 9820
rect 10909 9760 10973 9764
rect 10989 9820 11053 9824
rect 10989 9764 10993 9820
rect 10993 9764 11049 9820
rect 11049 9764 11053 9820
rect 10989 9760 11053 9764
rect 15648 9820 15712 9824
rect 15648 9764 15652 9820
rect 15652 9764 15708 9820
rect 15708 9764 15712 9820
rect 15648 9760 15712 9764
rect 15728 9820 15792 9824
rect 15728 9764 15732 9820
rect 15732 9764 15788 9820
rect 15788 9764 15792 9820
rect 15728 9760 15792 9764
rect 15808 9820 15872 9824
rect 15808 9764 15812 9820
rect 15812 9764 15868 9820
rect 15868 9764 15872 9820
rect 15808 9760 15872 9764
rect 15888 9820 15952 9824
rect 15888 9764 15892 9820
rect 15892 9764 15948 9820
rect 15948 9764 15952 9820
rect 15888 9760 15952 9764
rect 20547 9820 20611 9824
rect 20547 9764 20551 9820
rect 20551 9764 20607 9820
rect 20607 9764 20611 9820
rect 20547 9760 20611 9764
rect 20627 9820 20691 9824
rect 20627 9764 20631 9820
rect 20631 9764 20687 9820
rect 20687 9764 20691 9820
rect 20627 9760 20691 9764
rect 20707 9820 20771 9824
rect 20707 9764 20711 9820
rect 20711 9764 20767 9820
rect 20767 9764 20771 9820
rect 20707 9760 20771 9764
rect 20787 9820 20851 9824
rect 20787 9764 20791 9820
rect 20791 9764 20847 9820
rect 20847 9764 20851 9820
rect 20787 9760 20851 9764
rect 3401 9276 3465 9280
rect 3401 9220 3405 9276
rect 3405 9220 3461 9276
rect 3461 9220 3465 9276
rect 3401 9216 3465 9220
rect 3481 9276 3545 9280
rect 3481 9220 3485 9276
rect 3485 9220 3541 9276
rect 3541 9220 3545 9276
rect 3481 9216 3545 9220
rect 3561 9276 3625 9280
rect 3561 9220 3565 9276
rect 3565 9220 3621 9276
rect 3621 9220 3625 9276
rect 3561 9216 3625 9220
rect 3641 9276 3705 9280
rect 3641 9220 3645 9276
rect 3645 9220 3701 9276
rect 3701 9220 3705 9276
rect 3641 9216 3705 9220
rect 8300 9276 8364 9280
rect 8300 9220 8304 9276
rect 8304 9220 8360 9276
rect 8360 9220 8364 9276
rect 8300 9216 8364 9220
rect 8380 9276 8444 9280
rect 8380 9220 8384 9276
rect 8384 9220 8440 9276
rect 8440 9220 8444 9276
rect 8380 9216 8444 9220
rect 8460 9276 8524 9280
rect 8460 9220 8464 9276
rect 8464 9220 8520 9276
rect 8520 9220 8524 9276
rect 8460 9216 8524 9220
rect 8540 9276 8604 9280
rect 8540 9220 8544 9276
rect 8544 9220 8600 9276
rect 8600 9220 8604 9276
rect 8540 9216 8604 9220
rect 13199 9276 13263 9280
rect 13199 9220 13203 9276
rect 13203 9220 13259 9276
rect 13259 9220 13263 9276
rect 13199 9216 13263 9220
rect 13279 9276 13343 9280
rect 13279 9220 13283 9276
rect 13283 9220 13339 9276
rect 13339 9220 13343 9276
rect 13279 9216 13343 9220
rect 13359 9276 13423 9280
rect 13359 9220 13363 9276
rect 13363 9220 13419 9276
rect 13419 9220 13423 9276
rect 13359 9216 13423 9220
rect 13439 9276 13503 9280
rect 13439 9220 13443 9276
rect 13443 9220 13499 9276
rect 13499 9220 13503 9276
rect 13439 9216 13503 9220
rect 18098 9276 18162 9280
rect 18098 9220 18102 9276
rect 18102 9220 18158 9276
rect 18158 9220 18162 9276
rect 18098 9216 18162 9220
rect 18178 9276 18242 9280
rect 18178 9220 18182 9276
rect 18182 9220 18238 9276
rect 18238 9220 18242 9276
rect 18178 9216 18242 9220
rect 18258 9276 18322 9280
rect 18258 9220 18262 9276
rect 18262 9220 18318 9276
rect 18318 9220 18322 9276
rect 18258 9216 18322 9220
rect 18338 9276 18402 9280
rect 18338 9220 18342 9276
rect 18342 9220 18398 9276
rect 18398 9220 18402 9276
rect 18338 9216 18402 9220
rect 5850 8732 5914 8736
rect 5850 8676 5854 8732
rect 5854 8676 5910 8732
rect 5910 8676 5914 8732
rect 5850 8672 5914 8676
rect 5930 8732 5994 8736
rect 5930 8676 5934 8732
rect 5934 8676 5990 8732
rect 5990 8676 5994 8732
rect 5930 8672 5994 8676
rect 6010 8732 6074 8736
rect 6010 8676 6014 8732
rect 6014 8676 6070 8732
rect 6070 8676 6074 8732
rect 6010 8672 6074 8676
rect 6090 8732 6154 8736
rect 6090 8676 6094 8732
rect 6094 8676 6150 8732
rect 6150 8676 6154 8732
rect 6090 8672 6154 8676
rect 10749 8732 10813 8736
rect 10749 8676 10753 8732
rect 10753 8676 10809 8732
rect 10809 8676 10813 8732
rect 10749 8672 10813 8676
rect 10829 8732 10893 8736
rect 10829 8676 10833 8732
rect 10833 8676 10889 8732
rect 10889 8676 10893 8732
rect 10829 8672 10893 8676
rect 10909 8732 10973 8736
rect 10909 8676 10913 8732
rect 10913 8676 10969 8732
rect 10969 8676 10973 8732
rect 10909 8672 10973 8676
rect 10989 8732 11053 8736
rect 10989 8676 10993 8732
rect 10993 8676 11049 8732
rect 11049 8676 11053 8732
rect 10989 8672 11053 8676
rect 15648 8732 15712 8736
rect 15648 8676 15652 8732
rect 15652 8676 15708 8732
rect 15708 8676 15712 8732
rect 15648 8672 15712 8676
rect 15728 8732 15792 8736
rect 15728 8676 15732 8732
rect 15732 8676 15788 8732
rect 15788 8676 15792 8732
rect 15728 8672 15792 8676
rect 15808 8732 15872 8736
rect 15808 8676 15812 8732
rect 15812 8676 15868 8732
rect 15868 8676 15872 8732
rect 15808 8672 15872 8676
rect 15888 8732 15952 8736
rect 15888 8676 15892 8732
rect 15892 8676 15948 8732
rect 15948 8676 15952 8732
rect 15888 8672 15952 8676
rect 20547 8732 20611 8736
rect 20547 8676 20551 8732
rect 20551 8676 20607 8732
rect 20607 8676 20611 8732
rect 20547 8672 20611 8676
rect 20627 8732 20691 8736
rect 20627 8676 20631 8732
rect 20631 8676 20687 8732
rect 20687 8676 20691 8732
rect 20627 8672 20691 8676
rect 20707 8732 20771 8736
rect 20707 8676 20711 8732
rect 20711 8676 20767 8732
rect 20767 8676 20771 8732
rect 20707 8672 20771 8676
rect 20787 8732 20851 8736
rect 20787 8676 20791 8732
rect 20791 8676 20847 8732
rect 20847 8676 20851 8732
rect 20787 8672 20851 8676
rect 3401 8188 3465 8192
rect 3401 8132 3405 8188
rect 3405 8132 3461 8188
rect 3461 8132 3465 8188
rect 3401 8128 3465 8132
rect 3481 8188 3545 8192
rect 3481 8132 3485 8188
rect 3485 8132 3541 8188
rect 3541 8132 3545 8188
rect 3481 8128 3545 8132
rect 3561 8188 3625 8192
rect 3561 8132 3565 8188
rect 3565 8132 3621 8188
rect 3621 8132 3625 8188
rect 3561 8128 3625 8132
rect 3641 8188 3705 8192
rect 3641 8132 3645 8188
rect 3645 8132 3701 8188
rect 3701 8132 3705 8188
rect 3641 8128 3705 8132
rect 8300 8188 8364 8192
rect 8300 8132 8304 8188
rect 8304 8132 8360 8188
rect 8360 8132 8364 8188
rect 8300 8128 8364 8132
rect 8380 8188 8444 8192
rect 8380 8132 8384 8188
rect 8384 8132 8440 8188
rect 8440 8132 8444 8188
rect 8380 8128 8444 8132
rect 8460 8188 8524 8192
rect 8460 8132 8464 8188
rect 8464 8132 8520 8188
rect 8520 8132 8524 8188
rect 8460 8128 8524 8132
rect 8540 8188 8604 8192
rect 8540 8132 8544 8188
rect 8544 8132 8600 8188
rect 8600 8132 8604 8188
rect 8540 8128 8604 8132
rect 13199 8188 13263 8192
rect 13199 8132 13203 8188
rect 13203 8132 13259 8188
rect 13259 8132 13263 8188
rect 13199 8128 13263 8132
rect 13279 8188 13343 8192
rect 13279 8132 13283 8188
rect 13283 8132 13339 8188
rect 13339 8132 13343 8188
rect 13279 8128 13343 8132
rect 13359 8188 13423 8192
rect 13359 8132 13363 8188
rect 13363 8132 13419 8188
rect 13419 8132 13423 8188
rect 13359 8128 13423 8132
rect 13439 8188 13503 8192
rect 13439 8132 13443 8188
rect 13443 8132 13499 8188
rect 13499 8132 13503 8188
rect 13439 8128 13503 8132
rect 18098 8188 18162 8192
rect 18098 8132 18102 8188
rect 18102 8132 18158 8188
rect 18158 8132 18162 8188
rect 18098 8128 18162 8132
rect 18178 8188 18242 8192
rect 18178 8132 18182 8188
rect 18182 8132 18238 8188
rect 18238 8132 18242 8188
rect 18178 8128 18242 8132
rect 18258 8188 18322 8192
rect 18258 8132 18262 8188
rect 18262 8132 18318 8188
rect 18318 8132 18322 8188
rect 18258 8128 18322 8132
rect 18338 8188 18402 8192
rect 18338 8132 18342 8188
rect 18342 8132 18398 8188
rect 18398 8132 18402 8188
rect 18338 8128 18402 8132
rect 5850 7644 5914 7648
rect 5850 7588 5854 7644
rect 5854 7588 5910 7644
rect 5910 7588 5914 7644
rect 5850 7584 5914 7588
rect 5930 7644 5994 7648
rect 5930 7588 5934 7644
rect 5934 7588 5990 7644
rect 5990 7588 5994 7644
rect 5930 7584 5994 7588
rect 6010 7644 6074 7648
rect 6010 7588 6014 7644
rect 6014 7588 6070 7644
rect 6070 7588 6074 7644
rect 6010 7584 6074 7588
rect 6090 7644 6154 7648
rect 6090 7588 6094 7644
rect 6094 7588 6150 7644
rect 6150 7588 6154 7644
rect 6090 7584 6154 7588
rect 10749 7644 10813 7648
rect 10749 7588 10753 7644
rect 10753 7588 10809 7644
rect 10809 7588 10813 7644
rect 10749 7584 10813 7588
rect 10829 7644 10893 7648
rect 10829 7588 10833 7644
rect 10833 7588 10889 7644
rect 10889 7588 10893 7644
rect 10829 7584 10893 7588
rect 10909 7644 10973 7648
rect 10909 7588 10913 7644
rect 10913 7588 10969 7644
rect 10969 7588 10973 7644
rect 10909 7584 10973 7588
rect 10989 7644 11053 7648
rect 10989 7588 10993 7644
rect 10993 7588 11049 7644
rect 11049 7588 11053 7644
rect 10989 7584 11053 7588
rect 15648 7644 15712 7648
rect 15648 7588 15652 7644
rect 15652 7588 15708 7644
rect 15708 7588 15712 7644
rect 15648 7584 15712 7588
rect 15728 7644 15792 7648
rect 15728 7588 15732 7644
rect 15732 7588 15788 7644
rect 15788 7588 15792 7644
rect 15728 7584 15792 7588
rect 15808 7644 15872 7648
rect 15808 7588 15812 7644
rect 15812 7588 15868 7644
rect 15868 7588 15872 7644
rect 15808 7584 15872 7588
rect 15888 7644 15952 7648
rect 15888 7588 15892 7644
rect 15892 7588 15948 7644
rect 15948 7588 15952 7644
rect 15888 7584 15952 7588
rect 20547 7644 20611 7648
rect 20547 7588 20551 7644
rect 20551 7588 20607 7644
rect 20607 7588 20611 7644
rect 20547 7584 20611 7588
rect 20627 7644 20691 7648
rect 20627 7588 20631 7644
rect 20631 7588 20687 7644
rect 20687 7588 20691 7644
rect 20627 7584 20691 7588
rect 20707 7644 20771 7648
rect 20707 7588 20711 7644
rect 20711 7588 20767 7644
rect 20767 7588 20771 7644
rect 20707 7584 20771 7588
rect 20787 7644 20851 7648
rect 20787 7588 20791 7644
rect 20791 7588 20847 7644
rect 20847 7588 20851 7644
rect 20787 7584 20851 7588
rect 3401 7100 3465 7104
rect 3401 7044 3405 7100
rect 3405 7044 3461 7100
rect 3461 7044 3465 7100
rect 3401 7040 3465 7044
rect 3481 7100 3545 7104
rect 3481 7044 3485 7100
rect 3485 7044 3541 7100
rect 3541 7044 3545 7100
rect 3481 7040 3545 7044
rect 3561 7100 3625 7104
rect 3561 7044 3565 7100
rect 3565 7044 3621 7100
rect 3621 7044 3625 7100
rect 3561 7040 3625 7044
rect 3641 7100 3705 7104
rect 3641 7044 3645 7100
rect 3645 7044 3701 7100
rect 3701 7044 3705 7100
rect 3641 7040 3705 7044
rect 8300 7100 8364 7104
rect 8300 7044 8304 7100
rect 8304 7044 8360 7100
rect 8360 7044 8364 7100
rect 8300 7040 8364 7044
rect 8380 7100 8444 7104
rect 8380 7044 8384 7100
rect 8384 7044 8440 7100
rect 8440 7044 8444 7100
rect 8380 7040 8444 7044
rect 8460 7100 8524 7104
rect 8460 7044 8464 7100
rect 8464 7044 8520 7100
rect 8520 7044 8524 7100
rect 8460 7040 8524 7044
rect 8540 7100 8604 7104
rect 8540 7044 8544 7100
rect 8544 7044 8600 7100
rect 8600 7044 8604 7100
rect 8540 7040 8604 7044
rect 13199 7100 13263 7104
rect 13199 7044 13203 7100
rect 13203 7044 13259 7100
rect 13259 7044 13263 7100
rect 13199 7040 13263 7044
rect 13279 7100 13343 7104
rect 13279 7044 13283 7100
rect 13283 7044 13339 7100
rect 13339 7044 13343 7100
rect 13279 7040 13343 7044
rect 13359 7100 13423 7104
rect 13359 7044 13363 7100
rect 13363 7044 13419 7100
rect 13419 7044 13423 7100
rect 13359 7040 13423 7044
rect 13439 7100 13503 7104
rect 13439 7044 13443 7100
rect 13443 7044 13499 7100
rect 13499 7044 13503 7100
rect 13439 7040 13503 7044
rect 18098 7100 18162 7104
rect 18098 7044 18102 7100
rect 18102 7044 18158 7100
rect 18158 7044 18162 7100
rect 18098 7040 18162 7044
rect 18178 7100 18242 7104
rect 18178 7044 18182 7100
rect 18182 7044 18238 7100
rect 18238 7044 18242 7100
rect 18178 7040 18242 7044
rect 18258 7100 18322 7104
rect 18258 7044 18262 7100
rect 18262 7044 18318 7100
rect 18318 7044 18322 7100
rect 18258 7040 18322 7044
rect 18338 7100 18402 7104
rect 18338 7044 18342 7100
rect 18342 7044 18398 7100
rect 18398 7044 18402 7100
rect 18338 7040 18402 7044
rect 5850 6556 5914 6560
rect 5850 6500 5854 6556
rect 5854 6500 5910 6556
rect 5910 6500 5914 6556
rect 5850 6496 5914 6500
rect 5930 6556 5994 6560
rect 5930 6500 5934 6556
rect 5934 6500 5990 6556
rect 5990 6500 5994 6556
rect 5930 6496 5994 6500
rect 6010 6556 6074 6560
rect 6010 6500 6014 6556
rect 6014 6500 6070 6556
rect 6070 6500 6074 6556
rect 6010 6496 6074 6500
rect 6090 6556 6154 6560
rect 6090 6500 6094 6556
rect 6094 6500 6150 6556
rect 6150 6500 6154 6556
rect 6090 6496 6154 6500
rect 10749 6556 10813 6560
rect 10749 6500 10753 6556
rect 10753 6500 10809 6556
rect 10809 6500 10813 6556
rect 10749 6496 10813 6500
rect 10829 6556 10893 6560
rect 10829 6500 10833 6556
rect 10833 6500 10889 6556
rect 10889 6500 10893 6556
rect 10829 6496 10893 6500
rect 10909 6556 10973 6560
rect 10909 6500 10913 6556
rect 10913 6500 10969 6556
rect 10969 6500 10973 6556
rect 10909 6496 10973 6500
rect 10989 6556 11053 6560
rect 10989 6500 10993 6556
rect 10993 6500 11049 6556
rect 11049 6500 11053 6556
rect 10989 6496 11053 6500
rect 15648 6556 15712 6560
rect 15648 6500 15652 6556
rect 15652 6500 15708 6556
rect 15708 6500 15712 6556
rect 15648 6496 15712 6500
rect 15728 6556 15792 6560
rect 15728 6500 15732 6556
rect 15732 6500 15788 6556
rect 15788 6500 15792 6556
rect 15728 6496 15792 6500
rect 15808 6556 15872 6560
rect 15808 6500 15812 6556
rect 15812 6500 15868 6556
rect 15868 6500 15872 6556
rect 15808 6496 15872 6500
rect 15888 6556 15952 6560
rect 15888 6500 15892 6556
rect 15892 6500 15948 6556
rect 15948 6500 15952 6556
rect 15888 6496 15952 6500
rect 20547 6556 20611 6560
rect 20547 6500 20551 6556
rect 20551 6500 20607 6556
rect 20607 6500 20611 6556
rect 20547 6496 20611 6500
rect 20627 6556 20691 6560
rect 20627 6500 20631 6556
rect 20631 6500 20687 6556
rect 20687 6500 20691 6556
rect 20627 6496 20691 6500
rect 20707 6556 20771 6560
rect 20707 6500 20711 6556
rect 20711 6500 20767 6556
rect 20767 6500 20771 6556
rect 20707 6496 20771 6500
rect 20787 6556 20851 6560
rect 20787 6500 20791 6556
rect 20791 6500 20847 6556
rect 20847 6500 20851 6556
rect 20787 6496 20851 6500
rect 3401 6012 3465 6016
rect 3401 5956 3405 6012
rect 3405 5956 3461 6012
rect 3461 5956 3465 6012
rect 3401 5952 3465 5956
rect 3481 6012 3545 6016
rect 3481 5956 3485 6012
rect 3485 5956 3541 6012
rect 3541 5956 3545 6012
rect 3481 5952 3545 5956
rect 3561 6012 3625 6016
rect 3561 5956 3565 6012
rect 3565 5956 3621 6012
rect 3621 5956 3625 6012
rect 3561 5952 3625 5956
rect 3641 6012 3705 6016
rect 3641 5956 3645 6012
rect 3645 5956 3701 6012
rect 3701 5956 3705 6012
rect 3641 5952 3705 5956
rect 8300 6012 8364 6016
rect 8300 5956 8304 6012
rect 8304 5956 8360 6012
rect 8360 5956 8364 6012
rect 8300 5952 8364 5956
rect 8380 6012 8444 6016
rect 8380 5956 8384 6012
rect 8384 5956 8440 6012
rect 8440 5956 8444 6012
rect 8380 5952 8444 5956
rect 8460 6012 8524 6016
rect 8460 5956 8464 6012
rect 8464 5956 8520 6012
rect 8520 5956 8524 6012
rect 8460 5952 8524 5956
rect 8540 6012 8604 6016
rect 8540 5956 8544 6012
rect 8544 5956 8600 6012
rect 8600 5956 8604 6012
rect 8540 5952 8604 5956
rect 13199 6012 13263 6016
rect 13199 5956 13203 6012
rect 13203 5956 13259 6012
rect 13259 5956 13263 6012
rect 13199 5952 13263 5956
rect 13279 6012 13343 6016
rect 13279 5956 13283 6012
rect 13283 5956 13339 6012
rect 13339 5956 13343 6012
rect 13279 5952 13343 5956
rect 13359 6012 13423 6016
rect 13359 5956 13363 6012
rect 13363 5956 13419 6012
rect 13419 5956 13423 6012
rect 13359 5952 13423 5956
rect 13439 6012 13503 6016
rect 13439 5956 13443 6012
rect 13443 5956 13499 6012
rect 13499 5956 13503 6012
rect 13439 5952 13503 5956
rect 18098 6012 18162 6016
rect 18098 5956 18102 6012
rect 18102 5956 18158 6012
rect 18158 5956 18162 6012
rect 18098 5952 18162 5956
rect 18178 6012 18242 6016
rect 18178 5956 18182 6012
rect 18182 5956 18238 6012
rect 18238 5956 18242 6012
rect 18178 5952 18242 5956
rect 18258 6012 18322 6016
rect 18258 5956 18262 6012
rect 18262 5956 18318 6012
rect 18318 5956 18322 6012
rect 18258 5952 18322 5956
rect 18338 6012 18402 6016
rect 18338 5956 18342 6012
rect 18342 5956 18398 6012
rect 18398 5956 18402 6012
rect 18338 5952 18402 5956
rect 5850 5468 5914 5472
rect 5850 5412 5854 5468
rect 5854 5412 5910 5468
rect 5910 5412 5914 5468
rect 5850 5408 5914 5412
rect 5930 5468 5994 5472
rect 5930 5412 5934 5468
rect 5934 5412 5990 5468
rect 5990 5412 5994 5468
rect 5930 5408 5994 5412
rect 6010 5468 6074 5472
rect 6010 5412 6014 5468
rect 6014 5412 6070 5468
rect 6070 5412 6074 5468
rect 6010 5408 6074 5412
rect 6090 5468 6154 5472
rect 6090 5412 6094 5468
rect 6094 5412 6150 5468
rect 6150 5412 6154 5468
rect 6090 5408 6154 5412
rect 10749 5468 10813 5472
rect 10749 5412 10753 5468
rect 10753 5412 10809 5468
rect 10809 5412 10813 5468
rect 10749 5408 10813 5412
rect 10829 5468 10893 5472
rect 10829 5412 10833 5468
rect 10833 5412 10889 5468
rect 10889 5412 10893 5468
rect 10829 5408 10893 5412
rect 10909 5468 10973 5472
rect 10909 5412 10913 5468
rect 10913 5412 10969 5468
rect 10969 5412 10973 5468
rect 10909 5408 10973 5412
rect 10989 5468 11053 5472
rect 10989 5412 10993 5468
rect 10993 5412 11049 5468
rect 11049 5412 11053 5468
rect 10989 5408 11053 5412
rect 15648 5468 15712 5472
rect 15648 5412 15652 5468
rect 15652 5412 15708 5468
rect 15708 5412 15712 5468
rect 15648 5408 15712 5412
rect 15728 5468 15792 5472
rect 15728 5412 15732 5468
rect 15732 5412 15788 5468
rect 15788 5412 15792 5468
rect 15728 5408 15792 5412
rect 15808 5468 15872 5472
rect 15808 5412 15812 5468
rect 15812 5412 15868 5468
rect 15868 5412 15872 5468
rect 15808 5408 15872 5412
rect 15888 5468 15952 5472
rect 15888 5412 15892 5468
rect 15892 5412 15948 5468
rect 15948 5412 15952 5468
rect 15888 5408 15952 5412
rect 20547 5468 20611 5472
rect 20547 5412 20551 5468
rect 20551 5412 20607 5468
rect 20607 5412 20611 5468
rect 20547 5408 20611 5412
rect 20627 5468 20691 5472
rect 20627 5412 20631 5468
rect 20631 5412 20687 5468
rect 20687 5412 20691 5468
rect 20627 5408 20691 5412
rect 20707 5468 20771 5472
rect 20707 5412 20711 5468
rect 20711 5412 20767 5468
rect 20767 5412 20771 5468
rect 20707 5408 20771 5412
rect 20787 5468 20851 5472
rect 20787 5412 20791 5468
rect 20791 5412 20847 5468
rect 20847 5412 20851 5468
rect 20787 5408 20851 5412
rect 3401 4924 3465 4928
rect 3401 4868 3405 4924
rect 3405 4868 3461 4924
rect 3461 4868 3465 4924
rect 3401 4864 3465 4868
rect 3481 4924 3545 4928
rect 3481 4868 3485 4924
rect 3485 4868 3541 4924
rect 3541 4868 3545 4924
rect 3481 4864 3545 4868
rect 3561 4924 3625 4928
rect 3561 4868 3565 4924
rect 3565 4868 3621 4924
rect 3621 4868 3625 4924
rect 3561 4864 3625 4868
rect 3641 4924 3705 4928
rect 3641 4868 3645 4924
rect 3645 4868 3701 4924
rect 3701 4868 3705 4924
rect 3641 4864 3705 4868
rect 8300 4924 8364 4928
rect 8300 4868 8304 4924
rect 8304 4868 8360 4924
rect 8360 4868 8364 4924
rect 8300 4864 8364 4868
rect 8380 4924 8444 4928
rect 8380 4868 8384 4924
rect 8384 4868 8440 4924
rect 8440 4868 8444 4924
rect 8380 4864 8444 4868
rect 8460 4924 8524 4928
rect 8460 4868 8464 4924
rect 8464 4868 8520 4924
rect 8520 4868 8524 4924
rect 8460 4864 8524 4868
rect 8540 4924 8604 4928
rect 8540 4868 8544 4924
rect 8544 4868 8600 4924
rect 8600 4868 8604 4924
rect 8540 4864 8604 4868
rect 13199 4924 13263 4928
rect 13199 4868 13203 4924
rect 13203 4868 13259 4924
rect 13259 4868 13263 4924
rect 13199 4864 13263 4868
rect 13279 4924 13343 4928
rect 13279 4868 13283 4924
rect 13283 4868 13339 4924
rect 13339 4868 13343 4924
rect 13279 4864 13343 4868
rect 13359 4924 13423 4928
rect 13359 4868 13363 4924
rect 13363 4868 13419 4924
rect 13419 4868 13423 4924
rect 13359 4864 13423 4868
rect 13439 4924 13503 4928
rect 13439 4868 13443 4924
rect 13443 4868 13499 4924
rect 13499 4868 13503 4924
rect 13439 4864 13503 4868
rect 18098 4924 18162 4928
rect 18098 4868 18102 4924
rect 18102 4868 18158 4924
rect 18158 4868 18162 4924
rect 18098 4864 18162 4868
rect 18178 4924 18242 4928
rect 18178 4868 18182 4924
rect 18182 4868 18238 4924
rect 18238 4868 18242 4924
rect 18178 4864 18242 4868
rect 18258 4924 18322 4928
rect 18258 4868 18262 4924
rect 18262 4868 18318 4924
rect 18318 4868 18322 4924
rect 18258 4864 18322 4868
rect 18338 4924 18402 4928
rect 18338 4868 18342 4924
rect 18342 4868 18398 4924
rect 18398 4868 18402 4924
rect 18338 4864 18402 4868
rect 5850 4380 5914 4384
rect 5850 4324 5854 4380
rect 5854 4324 5910 4380
rect 5910 4324 5914 4380
rect 5850 4320 5914 4324
rect 5930 4380 5994 4384
rect 5930 4324 5934 4380
rect 5934 4324 5990 4380
rect 5990 4324 5994 4380
rect 5930 4320 5994 4324
rect 6010 4380 6074 4384
rect 6010 4324 6014 4380
rect 6014 4324 6070 4380
rect 6070 4324 6074 4380
rect 6010 4320 6074 4324
rect 6090 4380 6154 4384
rect 6090 4324 6094 4380
rect 6094 4324 6150 4380
rect 6150 4324 6154 4380
rect 6090 4320 6154 4324
rect 10749 4380 10813 4384
rect 10749 4324 10753 4380
rect 10753 4324 10809 4380
rect 10809 4324 10813 4380
rect 10749 4320 10813 4324
rect 10829 4380 10893 4384
rect 10829 4324 10833 4380
rect 10833 4324 10889 4380
rect 10889 4324 10893 4380
rect 10829 4320 10893 4324
rect 10909 4380 10973 4384
rect 10909 4324 10913 4380
rect 10913 4324 10969 4380
rect 10969 4324 10973 4380
rect 10909 4320 10973 4324
rect 10989 4380 11053 4384
rect 10989 4324 10993 4380
rect 10993 4324 11049 4380
rect 11049 4324 11053 4380
rect 10989 4320 11053 4324
rect 15648 4380 15712 4384
rect 15648 4324 15652 4380
rect 15652 4324 15708 4380
rect 15708 4324 15712 4380
rect 15648 4320 15712 4324
rect 15728 4380 15792 4384
rect 15728 4324 15732 4380
rect 15732 4324 15788 4380
rect 15788 4324 15792 4380
rect 15728 4320 15792 4324
rect 15808 4380 15872 4384
rect 15808 4324 15812 4380
rect 15812 4324 15868 4380
rect 15868 4324 15872 4380
rect 15808 4320 15872 4324
rect 15888 4380 15952 4384
rect 15888 4324 15892 4380
rect 15892 4324 15948 4380
rect 15948 4324 15952 4380
rect 15888 4320 15952 4324
rect 20547 4380 20611 4384
rect 20547 4324 20551 4380
rect 20551 4324 20607 4380
rect 20607 4324 20611 4380
rect 20547 4320 20611 4324
rect 20627 4380 20691 4384
rect 20627 4324 20631 4380
rect 20631 4324 20687 4380
rect 20687 4324 20691 4380
rect 20627 4320 20691 4324
rect 20707 4380 20771 4384
rect 20707 4324 20711 4380
rect 20711 4324 20767 4380
rect 20767 4324 20771 4380
rect 20707 4320 20771 4324
rect 20787 4380 20851 4384
rect 20787 4324 20791 4380
rect 20791 4324 20847 4380
rect 20847 4324 20851 4380
rect 20787 4320 20851 4324
rect 3401 3836 3465 3840
rect 3401 3780 3405 3836
rect 3405 3780 3461 3836
rect 3461 3780 3465 3836
rect 3401 3776 3465 3780
rect 3481 3836 3545 3840
rect 3481 3780 3485 3836
rect 3485 3780 3541 3836
rect 3541 3780 3545 3836
rect 3481 3776 3545 3780
rect 3561 3836 3625 3840
rect 3561 3780 3565 3836
rect 3565 3780 3621 3836
rect 3621 3780 3625 3836
rect 3561 3776 3625 3780
rect 3641 3836 3705 3840
rect 3641 3780 3645 3836
rect 3645 3780 3701 3836
rect 3701 3780 3705 3836
rect 3641 3776 3705 3780
rect 8300 3836 8364 3840
rect 8300 3780 8304 3836
rect 8304 3780 8360 3836
rect 8360 3780 8364 3836
rect 8300 3776 8364 3780
rect 8380 3836 8444 3840
rect 8380 3780 8384 3836
rect 8384 3780 8440 3836
rect 8440 3780 8444 3836
rect 8380 3776 8444 3780
rect 8460 3836 8524 3840
rect 8460 3780 8464 3836
rect 8464 3780 8520 3836
rect 8520 3780 8524 3836
rect 8460 3776 8524 3780
rect 8540 3836 8604 3840
rect 8540 3780 8544 3836
rect 8544 3780 8600 3836
rect 8600 3780 8604 3836
rect 8540 3776 8604 3780
rect 13199 3836 13263 3840
rect 13199 3780 13203 3836
rect 13203 3780 13259 3836
rect 13259 3780 13263 3836
rect 13199 3776 13263 3780
rect 13279 3836 13343 3840
rect 13279 3780 13283 3836
rect 13283 3780 13339 3836
rect 13339 3780 13343 3836
rect 13279 3776 13343 3780
rect 13359 3836 13423 3840
rect 13359 3780 13363 3836
rect 13363 3780 13419 3836
rect 13419 3780 13423 3836
rect 13359 3776 13423 3780
rect 13439 3836 13503 3840
rect 13439 3780 13443 3836
rect 13443 3780 13499 3836
rect 13499 3780 13503 3836
rect 13439 3776 13503 3780
rect 18098 3836 18162 3840
rect 18098 3780 18102 3836
rect 18102 3780 18158 3836
rect 18158 3780 18162 3836
rect 18098 3776 18162 3780
rect 18178 3836 18242 3840
rect 18178 3780 18182 3836
rect 18182 3780 18238 3836
rect 18238 3780 18242 3836
rect 18178 3776 18242 3780
rect 18258 3836 18322 3840
rect 18258 3780 18262 3836
rect 18262 3780 18318 3836
rect 18318 3780 18322 3836
rect 18258 3776 18322 3780
rect 18338 3836 18402 3840
rect 18338 3780 18342 3836
rect 18342 3780 18398 3836
rect 18398 3780 18402 3836
rect 18338 3776 18402 3780
rect 21220 3436 21284 3500
rect 5850 3292 5914 3296
rect 5850 3236 5854 3292
rect 5854 3236 5910 3292
rect 5910 3236 5914 3292
rect 5850 3232 5914 3236
rect 5930 3292 5994 3296
rect 5930 3236 5934 3292
rect 5934 3236 5990 3292
rect 5990 3236 5994 3292
rect 5930 3232 5994 3236
rect 6010 3292 6074 3296
rect 6010 3236 6014 3292
rect 6014 3236 6070 3292
rect 6070 3236 6074 3292
rect 6010 3232 6074 3236
rect 6090 3292 6154 3296
rect 6090 3236 6094 3292
rect 6094 3236 6150 3292
rect 6150 3236 6154 3292
rect 6090 3232 6154 3236
rect 10749 3292 10813 3296
rect 10749 3236 10753 3292
rect 10753 3236 10809 3292
rect 10809 3236 10813 3292
rect 10749 3232 10813 3236
rect 10829 3292 10893 3296
rect 10829 3236 10833 3292
rect 10833 3236 10889 3292
rect 10889 3236 10893 3292
rect 10829 3232 10893 3236
rect 10909 3292 10973 3296
rect 10909 3236 10913 3292
rect 10913 3236 10969 3292
rect 10969 3236 10973 3292
rect 10909 3232 10973 3236
rect 10989 3292 11053 3296
rect 10989 3236 10993 3292
rect 10993 3236 11049 3292
rect 11049 3236 11053 3292
rect 10989 3232 11053 3236
rect 15648 3292 15712 3296
rect 15648 3236 15652 3292
rect 15652 3236 15708 3292
rect 15708 3236 15712 3292
rect 15648 3232 15712 3236
rect 15728 3292 15792 3296
rect 15728 3236 15732 3292
rect 15732 3236 15788 3292
rect 15788 3236 15792 3292
rect 15728 3232 15792 3236
rect 15808 3292 15872 3296
rect 15808 3236 15812 3292
rect 15812 3236 15868 3292
rect 15868 3236 15872 3292
rect 15808 3232 15872 3236
rect 15888 3292 15952 3296
rect 15888 3236 15892 3292
rect 15892 3236 15948 3292
rect 15948 3236 15952 3292
rect 15888 3232 15952 3236
rect 20547 3292 20611 3296
rect 20547 3236 20551 3292
rect 20551 3236 20607 3292
rect 20607 3236 20611 3292
rect 20547 3232 20611 3236
rect 20627 3292 20691 3296
rect 20627 3236 20631 3292
rect 20631 3236 20687 3292
rect 20687 3236 20691 3292
rect 20627 3232 20691 3236
rect 20707 3292 20771 3296
rect 20707 3236 20711 3292
rect 20711 3236 20767 3292
rect 20767 3236 20771 3292
rect 20707 3232 20771 3236
rect 20787 3292 20851 3296
rect 20787 3236 20791 3292
rect 20791 3236 20847 3292
rect 20847 3236 20851 3292
rect 20787 3232 20851 3236
rect 21220 3164 21284 3228
rect 3401 2748 3465 2752
rect 3401 2692 3405 2748
rect 3405 2692 3461 2748
rect 3461 2692 3465 2748
rect 3401 2688 3465 2692
rect 3481 2748 3545 2752
rect 3481 2692 3485 2748
rect 3485 2692 3541 2748
rect 3541 2692 3545 2748
rect 3481 2688 3545 2692
rect 3561 2748 3625 2752
rect 3561 2692 3565 2748
rect 3565 2692 3621 2748
rect 3621 2692 3625 2748
rect 3561 2688 3625 2692
rect 3641 2748 3705 2752
rect 3641 2692 3645 2748
rect 3645 2692 3701 2748
rect 3701 2692 3705 2748
rect 3641 2688 3705 2692
rect 8300 2748 8364 2752
rect 8300 2692 8304 2748
rect 8304 2692 8360 2748
rect 8360 2692 8364 2748
rect 8300 2688 8364 2692
rect 8380 2748 8444 2752
rect 8380 2692 8384 2748
rect 8384 2692 8440 2748
rect 8440 2692 8444 2748
rect 8380 2688 8444 2692
rect 8460 2748 8524 2752
rect 8460 2692 8464 2748
rect 8464 2692 8520 2748
rect 8520 2692 8524 2748
rect 8460 2688 8524 2692
rect 8540 2748 8604 2752
rect 8540 2692 8544 2748
rect 8544 2692 8600 2748
rect 8600 2692 8604 2748
rect 8540 2688 8604 2692
rect 13199 2748 13263 2752
rect 13199 2692 13203 2748
rect 13203 2692 13259 2748
rect 13259 2692 13263 2748
rect 13199 2688 13263 2692
rect 13279 2748 13343 2752
rect 13279 2692 13283 2748
rect 13283 2692 13339 2748
rect 13339 2692 13343 2748
rect 13279 2688 13343 2692
rect 13359 2748 13423 2752
rect 13359 2692 13363 2748
rect 13363 2692 13419 2748
rect 13419 2692 13423 2748
rect 13359 2688 13423 2692
rect 13439 2748 13503 2752
rect 13439 2692 13443 2748
rect 13443 2692 13499 2748
rect 13499 2692 13503 2748
rect 13439 2688 13503 2692
rect 18098 2748 18162 2752
rect 18098 2692 18102 2748
rect 18102 2692 18158 2748
rect 18158 2692 18162 2748
rect 18098 2688 18162 2692
rect 18178 2748 18242 2752
rect 18178 2692 18182 2748
rect 18182 2692 18238 2748
rect 18238 2692 18242 2748
rect 18178 2688 18242 2692
rect 18258 2748 18322 2752
rect 18258 2692 18262 2748
rect 18262 2692 18318 2748
rect 18318 2692 18322 2748
rect 18258 2688 18322 2692
rect 18338 2748 18402 2752
rect 18338 2692 18342 2748
rect 18342 2692 18398 2748
rect 18398 2692 18402 2748
rect 18338 2688 18402 2692
rect 5850 2204 5914 2208
rect 5850 2148 5854 2204
rect 5854 2148 5910 2204
rect 5910 2148 5914 2204
rect 5850 2144 5914 2148
rect 5930 2204 5994 2208
rect 5930 2148 5934 2204
rect 5934 2148 5990 2204
rect 5990 2148 5994 2204
rect 5930 2144 5994 2148
rect 6010 2204 6074 2208
rect 6010 2148 6014 2204
rect 6014 2148 6070 2204
rect 6070 2148 6074 2204
rect 6010 2144 6074 2148
rect 6090 2204 6154 2208
rect 6090 2148 6094 2204
rect 6094 2148 6150 2204
rect 6150 2148 6154 2204
rect 6090 2144 6154 2148
rect 10749 2204 10813 2208
rect 10749 2148 10753 2204
rect 10753 2148 10809 2204
rect 10809 2148 10813 2204
rect 10749 2144 10813 2148
rect 10829 2204 10893 2208
rect 10829 2148 10833 2204
rect 10833 2148 10889 2204
rect 10889 2148 10893 2204
rect 10829 2144 10893 2148
rect 10909 2204 10973 2208
rect 10909 2148 10913 2204
rect 10913 2148 10969 2204
rect 10969 2148 10973 2204
rect 10909 2144 10973 2148
rect 10989 2204 11053 2208
rect 10989 2148 10993 2204
rect 10993 2148 11049 2204
rect 11049 2148 11053 2204
rect 10989 2144 11053 2148
rect 15648 2204 15712 2208
rect 15648 2148 15652 2204
rect 15652 2148 15708 2204
rect 15708 2148 15712 2204
rect 15648 2144 15712 2148
rect 15728 2204 15792 2208
rect 15728 2148 15732 2204
rect 15732 2148 15788 2204
rect 15788 2148 15792 2204
rect 15728 2144 15792 2148
rect 15808 2204 15872 2208
rect 15808 2148 15812 2204
rect 15812 2148 15868 2204
rect 15868 2148 15872 2204
rect 15808 2144 15872 2148
rect 15888 2204 15952 2208
rect 15888 2148 15892 2204
rect 15892 2148 15948 2204
rect 15948 2148 15952 2204
rect 15888 2144 15952 2148
rect 20547 2204 20611 2208
rect 20547 2148 20551 2204
rect 20551 2148 20607 2204
rect 20607 2148 20611 2204
rect 20547 2144 20611 2148
rect 20627 2204 20691 2208
rect 20627 2148 20631 2204
rect 20631 2148 20687 2204
rect 20687 2148 20691 2204
rect 20627 2144 20691 2148
rect 20707 2204 20771 2208
rect 20707 2148 20711 2204
rect 20711 2148 20767 2204
rect 20767 2148 20771 2204
rect 20707 2144 20771 2148
rect 20787 2204 20851 2208
rect 20787 2148 20791 2204
rect 20791 2148 20847 2204
rect 20847 2148 20851 2204
rect 20787 2144 20851 2148
<< metal4 >>
rect 3393 21248 3713 21808
rect 3393 21184 3401 21248
rect 3465 21184 3481 21248
rect 3545 21184 3561 21248
rect 3625 21184 3641 21248
rect 3705 21184 3713 21248
rect 3393 20160 3713 21184
rect 3393 20096 3401 20160
rect 3465 20096 3481 20160
rect 3545 20096 3561 20160
rect 3625 20096 3641 20160
rect 3705 20096 3713 20160
rect 3393 19072 3713 20096
rect 3393 19008 3401 19072
rect 3465 19008 3481 19072
rect 3545 19008 3561 19072
rect 3625 19008 3641 19072
rect 3705 19008 3713 19072
rect 3393 17984 3713 19008
rect 3393 17920 3401 17984
rect 3465 17920 3481 17984
rect 3545 17920 3561 17984
rect 3625 17920 3641 17984
rect 3705 17920 3713 17984
rect 3393 16896 3713 17920
rect 3393 16832 3401 16896
rect 3465 16832 3481 16896
rect 3545 16832 3561 16896
rect 3625 16832 3641 16896
rect 3705 16832 3713 16896
rect 3393 15808 3713 16832
rect 3393 15744 3401 15808
rect 3465 15744 3481 15808
rect 3545 15744 3561 15808
rect 3625 15744 3641 15808
rect 3705 15744 3713 15808
rect 3393 14720 3713 15744
rect 3393 14656 3401 14720
rect 3465 14656 3481 14720
rect 3545 14656 3561 14720
rect 3625 14656 3641 14720
rect 3705 14656 3713 14720
rect 3393 13632 3713 14656
rect 3393 13568 3401 13632
rect 3465 13568 3481 13632
rect 3545 13568 3561 13632
rect 3625 13568 3641 13632
rect 3705 13568 3713 13632
rect 3393 12544 3713 13568
rect 3393 12480 3401 12544
rect 3465 12480 3481 12544
rect 3545 12480 3561 12544
rect 3625 12480 3641 12544
rect 3705 12480 3713 12544
rect 3393 11456 3713 12480
rect 3393 11392 3401 11456
rect 3465 11392 3481 11456
rect 3545 11392 3561 11456
rect 3625 11392 3641 11456
rect 3705 11392 3713 11456
rect 3393 10368 3713 11392
rect 3393 10304 3401 10368
rect 3465 10304 3481 10368
rect 3545 10304 3561 10368
rect 3625 10304 3641 10368
rect 3705 10304 3713 10368
rect 3393 9280 3713 10304
rect 3393 9216 3401 9280
rect 3465 9216 3481 9280
rect 3545 9216 3561 9280
rect 3625 9216 3641 9280
rect 3705 9216 3713 9280
rect 3393 8192 3713 9216
rect 3393 8128 3401 8192
rect 3465 8128 3481 8192
rect 3545 8128 3561 8192
rect 3625 8128 3641 8192
rect 3705 8128 3713 8192
rect 3393 7104 3713 8128
rect 3393 7040 3401 7104
rect 3465 7040 3481 7104
rect 3545 7040 3561 7104
rect 3625 7040 3641 7104
rect 3705 7040 3713 7104
rect 3393 6016 3713 7040
rect 3393 5952 3401 6016
rect 3465 5952 3481 6016
rect 3545 5952 3561 6016
rect 3625 5952 3641 6016
rect 3705 5952 3713 6016
rect 3393 4928 3713 5952
rect 3393 4864 3401 4928
rect 3465 4864 3481 4928
rect 3545 4864 3561 4928
rect 3625 4864 3641 4928
rect 3705 4864 3713 4928
rect 3393 3840 3713 4864
rect 3393 3776 3401 3840
rect 3465 3776 3481 3840
rect 3545 3776 3561 3840
rect 3625 3776 3641 3840
rect 3705 3776 3713 3840
rect 3393 2752 3713 3776
rect 3393 2688 3401 2752
rect 3465 2688 3481 2752
rect 3545 2688 3561 2752
rect 3625 2688 3641 2752
rect 3705 2688 3713 2752
rect 3393 2128 3713 2688
rect 5842 21792 6162 21808
rect 5842 21728 5850 21792
rect 5914 21728 5930 21792
rect 5994 21728 6010 21792
rect 6074 21728 6090 21792
rect 6154 21728 6162 21792
rect 5842 20704 6162 21728
rect 5842 20640 5850 20704
rect 5914 20640 5930 20704
rect 5994 20640 6010 20704
rect 6074 20640 6090 20704
rect 6154 20640 6162 20704
rect 5842 19616 6162 20640
rect 5842 19552 5850 19616
rect 5914 19552 5930 19616
rect 5994 19552 6010 19616
rect 6074 19552 6090 19616
rect 6154 19552 6162 19616
rect 5842 18528 6162 19552
rect 5842 18464 5850 18528
rect 5914 18464 5930 18528
rect 5994 18464 6010 18528
rect 6074 18464 6090 18528
rect 6154 18464 6162 18528
rect 5842 17440 6162 18464
rect 5842 17376 5850 17440
rect 5914 17376 5930 17440
rect 5994 17376 6010 17440
rect 6074 17376 6090 17440
rect 6154 17376 6162 17440
rect 5842 16352 6162 17376
rect 5842 16288 5850 16352
rect 5914 16288 5930 16352
rect 5994 16288 6010 16352
rect 6074 16288 6090 16352
rect 6154 16288 6162 16352
rect 5842 15264 6162 16288
rect 5842 15200 5850 15264
rect 5914 15200 5930 15264
rect 5994 15200 6010 15264
rect 6074 15200 6090 15264
rect 6154 15200 6162 15264
rect 5842 14176 6162 15200
rect 5842 14112 5850 14176
rect 5914 14112 5930 14176
rect 5994 14112 6010 14176
rect 6074 14112 6090 14176
rect 6154 14112 6162 14176
rect 5842 13088 6162 14112
rect 5842 13024 5850 13088
rect 5914 13024 5930 13088
rect 5994 13024 6010 13088
rect 6074 13024 6090 13088
rect 6154 13024 6162 13088
rect 5842 12000 6162 13024
rect 5842 11936 5850 12000
rect 5914 11936 5930 12000
rect 5994 11936 6010 12000
rect 6074 11936 6090 12000
rect 6154 11936 6162 12000
rect 5842 10912 6162 11936
rect 5842 10848 5850 10912
rect 5914 10848 5930 10912
rect 5994 10848 6010 10912
rect 6074 10848 6090 10912
rect 6154 10848 6162 10912
rect 5842 9824 6162 10848
rect 5842 9760 5850 9824
rect 5914 9760 5930 9824
rect 5994 9760 6010 9824
rect 6074 9760 6090 9824
rect 6154 9760 6162 9824
rect 5842 8736 6162 9760
rect 5842 8672 5850 8736
rect 5914 8672 5930 8736
rect 5994 8672 6010 8736
rect 6074 8672 6090 8736
rect 6154 8672 6162 8736
rect 5842 7648 6162 8672
rect 5842 7584 5850 7648
rect 5914 7584 5930 7648
rect 5994 7584 6010 7648
rect 6074 7584 6090 7648
rect 6154 7584 6162 7648
rect 5842 6560 6162 7584
rect 5842 6496 5850 6560
rect 5914 6496 5930 6560
rect 5994 6496 6010 6560
rect 6074 6496 6090 6560
rect 6154 6496 6162 6560
rect 5842 5472 6162 6496
rect 5842 5408 5850 5472
rect 5914 5408 5930 5472
rect 5994 5408 6010 5472
rect 6074 5408 6090 5472
rect 6154 5408 6162 5472
rect 5842 4384 6162 5408
rect 5842 4320 5850 4384
rect 5914 4320 5930 4384
rect 5994 4320 6010 4384
rect 6074 4320 6090 4384
rect 6154 4320 6162 4384
rect 5842 3296 6162 4320
rect 5842 3232 5850 3296
rect 5914 3232 5930 3296
rect 5994 3232 6010 3296
rect 6074 3232 6090 3296
rect 6154 3232 6162 3296
rect 5842 2208 6162 3232
rect 5842 2144 5850 2208
rect 5914 2144 5930 2208
rect 5994 2144 6010 2208
rect 6074 2144 6090 2208
rect 6154 2144 6162 2208
rect 5842 2128 6162 2144
rect 8292 21248 8612 21808
rect 8292 21184 8300 21248
rect 8364 21184 8380 21248
rect 8444 21184 8460 21248
rect 8524 21184 8540 21248
rect 8604 21184 8612 21248
rect 8292 20160 8612 21184
rect 8292 20096 8300 20160
rect 8364 20096 8380 20160
rect 8444 20096 8460 20160
rect 8524 20096 8540 20160
rect 8604 20096 8612 20160
rect 8292 19072 8612 20096
rect 8292 19008 8300 19072
rect 8364 19008 8380 19072
rect 8444 19008 8460 19072
rect 8524 19008 8540 19072
rect 8604 19008 8612 19072
rect 8292 17984 8612 19008
rect 8292 17920 8300 17984
rect 8364 17920 8380 17984
rect 8444 17920 8460 17984
rect 8524 17920 8540 17984
rect 8604 17920 8612 17984
rect 8292 16896 8612 17920
rect 8292 16832 8300 16896
rect 8364 16832 8380 16896
rect 8444 16832 8460 16896
rect 8524 16832 8540 16896
rect 8604 16832 8612 16896
rect 8292 15808 8612 16832
rect 8292 15744 8300 15808
rect 8364 15744 8380 15808
rect 8444 15744 8460 15808
rect 8524 15744 8540 15808
rect 8604 15744 8612 15808
rect 8292 14720 8612 15744
rect 8292 14656 8300 14720
rect 8364 14656 8380 14720
rect 8444 14656 8460 14720
rect 8524 14656 8540 14720
rect 8604 14656 8612 14720
rect 8292 13632 8612 14656
rect 8292 13568 8300 13632
rect 8364 13568 8380 13632
rect 8444 13568 8460 13632
rect 8524 13568 8540 13632
rect 8604 13568 8612 13632
rect 8292 12544 8612 13568
rect 8292 12480 8300 12544
rect 8364 12480 8380 12544
rect 8444 12480 8460 12544
rect 8524 12480 8540 12544
rect 8604 12480 8612 12544
rect 8292 11456 8612 12480
rect 8292 11392 8300 11456
rect 8364 11392 8380 11456
rect 8444 11392 8460 11456
rect 8524 11392 8540 11456
rect 8604 11392 8612 11456
rect 8292 10368 8612 11392
rect 8292 10304 8300 10368
rect 8364 10304 8380 10368
rect 8444 10304 8460 10368
rect 8524 10304 8540 10368
rect 8604 10304 8612 10368
rect 8292 9280 8612 10304
rect 8292 9216 8300 9280
rect 8364 9216 8380 9280
rect 8444 9216 8460 9280
rect 8524 9216 8540 9280
rect 8604 9216 8612 9280
rect 8292 8192 8612 9216
rect 8292 8128 8300 8192
rect 8364 8128 8380 8192
rect 8444 8128 8460 8192
rect 8524 8128 8540 8192
rect 8604 8128 8612 8192
rect 8292 7104 8612 8128
rect 8292 7040 8300 7104
rect 8364 7040 8380 7104
rect 8444 7040 8460 7104
rect 8524 7040 8540 7104
rect 8604 7040 8612 7104
rect 8292 6016 8612 7040
rect 8292 5952 8300 6016
rect 8364 5952 8380 6016
rect 8444 5952 8460 6016
rect 8524 5952 8540 6016
rect 8604 5952 8612 6016
rect 8292 4928 8612 5952
rect 8292 4864 8300 4928
rect 8364 4864 8380 4928
rect 8444 4864 8460 4928
rect 8524 4864 8540 4928
rect 8604 4864 8612 4928
rect 8292 3840 8612 4864
rect 8292 3776 8300 3840
rect 8364 3776 8380 3840
rect 8444 3776 8460 3840
rect 8524 3776 8540 3840
rect 8604 3776 8612 3840
rect 8292 2752 8612 3776
rect 8292 2688 8300 2752
rect 8364 2688 8380 2752
rect 8444 2688 8460 2752
rect 8524 2688 8540 2752
rect 8604 2688 8612 2752
rect 8292 2128 8612 2688
rect 10741 21792 11061 21808
rect 10741 21728 10749 21792
rect 10813 21728 10829 21792
rect 10893 21728 10909 21792
rect 10973 21728 10989 21792
rect 11053 21728 11061 21792
rect 10741 20704 11061 21728
rect 10741 20640 10749 20704
rect 10813 20640 10829 20704
rect 10893 20640 10909 20704
rect 10973 20640 10989 20704
rect 11053 20640 11061 20704
rect 10741 19616 11061 20640
rect 10741 19552 10749 19616
rect 10813 19552 10829 19616
rect 10893 19552 10909 19616
rect 10973 19552 10989 19616
rect 11053 19552 11061 19616
rect 10741 18528 11061 19552
rect 10741 18464 10749 18528
rect 10813 18464 10829 18528
rect 10893 18464 10909 18528
rect 10973 18464 10989 18528
rect 11053 18464 11061 18528
rect 10741 17440 11061 18464
rect 10741 17376 10749 17440
rect 10813 17376 10829 17440
rect 10893 17376 10909 17440
rect 10973 17376 10989 17440
rect 11053 17376 11061 17440
rect 10741 16352 11061 17376
rect 10741 16288 10749 16352
rect 10813 16288 10829 16352
rect 10893 16288 10909 16352
rect 10973 16288 10989 16352
rect 11053 16288 11061 16352
rect 10741 15264 11061 16288
rect 10741 15200 10749 15264
rect 10813 15200 10829 15264
rect 10893 15200 10909 15264
rect 10973 15200 10989 15264
rect 11053 15200 11061 15264
rect 10741 14176 11061 15200
rect 10741 14112 10749 14176
rect 10813 14112 10829 14176
rect 10893 14112 10909 14176
rect 10973 14112 10989 14176
rect 11053 14112 11061 14176
rect 10741 13088 11061 14112
rect 10741 13024 10749 13088
rect 10813 13024 10829 13088
rect 10893 13024 10909 13088
rect 10973 13024 10989 13088
rect 11053 13024 11061 13088
rect 10741 12000 11061 13024
rect 10741 11936 10749 12000
rect 10813 11936 10829 12000
rect 10893 11936 10909 12000
rect 10973 11936 10989 12000
rect 11053 11936 11061 12000
rect 10741 10912 11061 11936
rect 10741 10848 10749 10912
rect 10813 10848 10829 10912
rect 10893 10848 10909 10912
rect 10973 10848 10989 10912
rect 11053 10848 11061 10912
rect 10741 9824 11061 10848
rect 10741 9760 10749 9824
rect 10813 9760 10829 9824
rect 10893 9760 10909 9824
rect 10973 9760 10989 9824
rect 11053 9760 11061 9824
rect 10741 8736 11061 9760
rect 10741 8672 10749 8736
rect 10813 8672 10829 8736
rect 10893 8672 10909 8736
rect 10973 8672 10989 8736
rect 11053 8672 11061 8736
rect 10741 7648 11061 8672
rect 10741 7584 10749 7648
rect 10813 7584 10829 7648
rect 10893 7584 10909 7648
rect 10973 7584 10989 7648
rect 11053 7584 11061 7648
rect 10741 6560 11061 7584
rect 10741 6496 10749 6560
rect 10813 6496 10829 6560
rect 10893 6496 10909 6560
rect 10973 6496 10989 6560
rect 11053 6496 11061 6560
rect 10741 5472 11061 6496
rect 10741 5408 10749 5472
rect 10813 5408 10829 5472
rect 10893 5408 10909 5472
rect 10973 5408 10989 5472
rect 11053 5408 11061 5472
rect 10741 4384 11061 5408
rect 10741 4320 10749 4384
rect 10813 4320 10829 4384
rect 10893 4320 10909 4384
rect 10973 4320 10989 4384
rect 11053 4320 11061 4384
rect 10741 3296 11061 4320
rect 10741 3232 10749 3296
rect 10813 3232 10829 3296
rect 10893 3232 10909 3296
rect 10973 3232 10989 3296
rect 11053 3232 11061 3296
rect 10741 2208 11061 3232
rect 10741 2144 10749 2208
rect 10813 2144 10829 2208
rect 10893 2144 10909 2208
rect 10973 2144 10989 2208
rect 11053 2144 11061 2208
rect 10741 2128 11061 2144
rect 13191 21248 13511 21808
rect 13191 21184 13199 21248
rect 13263 21184 13279 21248
rect 13343 21184 13359 21248
rect 13423 21184 13439 21248
rect 13503 21184 13511 21248
rect 13191 20160 13511 21184
rect 13191 20096 13199 20160
rect 13263 20096 13279 20160
rect 13343 20096 13359 20160
rect 13423 20096 13439 20160
rect 13503 20096 13511 20160
rect 13191 19072 13511 20096
rect 13191 19008 13199 19072
rect 13263 19008 13279 19072
rect 13343 19008 13359 19072
rect 13423 19008 13439 19072
rect 13503 19008 13511 19072
rect 13191 17984 13511 19008
rect 13191 17920 13199 17984
rect 13263 17920 13279 17984
rect 13343 17920 13359 17984
rect 13423 17920 13439 17984
rect 13503 17920 13511 17984
rect 13191 16896 13511 17920
rect 13191 16832 13199 16896
rect 13263 16832 13279 16896
rect 13343 16832 13359 16896
rect 13423 16832 13439 16896
rect 13503 16832 13511 16896
rect 13191 15808 13511 16832
rect 13191 15744 13199 15808
rect 13263 15744 13279 15808
rect 13343 15744 13359 15808
rect 13423 15744 13439 15808
rect 13503 15744 13511 15808
rect 13191 14720 13511 15744
rect 13191 14656 13199 14720
rect 13263 14656 13279 14720
rect 13343 14656 13359 14720
rect 13423 14656 13439 14720
rect 13503 14656 13511 14720
rect 13191 13632 13511 14656
rect 13191 13568 13199 13632
rect 13263 13568 13279 13632
rect 13343 13568 13359 13632
rect 13423 13568 13439 13632
rect 13503 13568 13511 13632
rect 13191 12544 13511 13568
rect 13191 12480 13199 12544
rect 13263 12480 13279 12544
rect 13343 12480 13359 12544
rect 13423 12480 13439 12544
rect 13503 12480 13511 12544
rect 13191 11456 13511 12480
rect 13191 11392 13199 11456
rect 13263 11392 13279 11456
rect 13343 11392 13359 11456
rect 13423 11392 13439 11456
rect 13503 11392 13511 11456
rect 13191 10368 13511 11392
rect 13191 10304 13199 10368
rect 13263 10304 13279 10368
rect 13343 10304 13359 10368
rect 13423 10304 13439 10368
rect 13503 10304 13511 10368
rect 13191 9280 13511 10304
rect 13191 9216 13199 9280
rect 13263 9216 13279 9280
rect 13343 9216 13359 9280
rect 13423 9216 13439 9280
rect 13503 9216 13511 9280
rect 13191 8192 13511 9216
rect 13191 8128 13199 8192
rect 13263 8128 13279 8192
rect 13343 8128 13359 8192
rect 13423 8128 13439 8192
rect 13503 8128 13511 8192
rect 13191 7104 13511 8128
rect 13191 7040 13199 7104
rect 13263 7040 13279 7104
rect 13343 7040 13359 7104
rect 13423 7040 13439 7104
rect 13503 7040 13511 7104
rect 13191 6016 13511 7040
rect 13191 5952 13199 6016
rect 13263 5952 13279 6016
rect 13343 5952 13359 6016
rect 13423 5952 13439 6016
rect 13503 5952 13511 6016
rect 13191 4928 13511 5952
rect 13191 4864 13199 4928
rect 13263 4864 13279 4928
rect 13343 4864 13359 4928
rect 13423 4864 13439 4928
rect 13503 4864 13511 4928
rect 13191 3840 13511 4864
rect 13191 3776 13199 3840
rect 13263 3776 13279 3840
rect 13343 3776 13359 3840
rect 13423 3776 13439 3840
rect 13503 3776 13511 3840
rect 13191 2752 13511 3776
rect 13191 2688 13199 2752
rect 13263 2688 13279 2752
rect 13343 2688 13359 2752
rect 13423 2688 13439 2752
rect 13503 2688 13511 2752
rect 13191 2128 13511 2688
rect 15640 21792 15960 21808
rect 15640 21728 15648 21792
rect 15712 21728 15728 21792
rect 15792 21728 15808 21792
rect 15872 21728 15888 21792
rect 15952 21728 15960 21792
rect 15640 20704 15960 21728
rect 15640 20640 15648 20704
rect 15712 20640 15728 20704
rect 15792 20640 15808 20704
rect 15872 20640 15888 20704
rect 15952 20640 15960 20704
rect 15640 19616 15960 20640
rect 15640 19552 15648 19616
rect 15712 19552 15728 19616
rect 15792 19552 15808 19616
rect 15872 19552 15888 19616
rect 15952 19552 15960 19616
rect 15640 18528 15960 19552
rect 15640 18464 15648 18528
rect 15712 18464 15728 18528
rect 15792 18464 15808 18528
rect 15872 18464 15888 18528
rect 15952 18464 15960 18528
rect 15640 17440 15960 18464
rect 15640 17376 15648 17440
rect 15712 17376 15728 17440
rect 15792 17376 15808 17440
rect 15872 17376 15888 17440
rect 15952 17376 15960 17440
rect 15640 16352 15960 17376
rect 15640 16288 15648 16352
rect 15712 16288 15728 16352
rect 15792 16288 15808 16352
rect 15872 16288 15888 16352
rect 15952 16288 15960 16352
rect 15640 15264 15960 16288
rect 15640 15200 15648 15264
rect 15712 15200 15728 15264
rect 15792 15200 15808 15264
rect 15872 15200 15888 15264
rect 15952 15200 15960 15264
rect 15640 14176 15960 15200
rect 15640 14112 15648 14176
rect 15712 14112 15728 14176
rect 15792 14112 15808 14176
rect 15872 14112 15888 14176
rect 15952 14112 15960 14176
rect 15640 13088 15960 14112
rect 15640 13024 15648 13088
rect 15712 13024 15728 13088
rect 15792 13024 15808 13088
rect 15872 13024 15888 13088
rect 15952 13024 15960 13088
rect 15640 12000 15960 13024
rect 15640 11936 15648 12000
rect 15712 11936 15728 12000
rect 15792 11936 15808 12000
rect 15872 11936 15888 12000
rect 15952 11936 15960 12000
rect 15640 10912 15960 11936
rect 15640 10848 15648 10912
rect 15712 10848 15728 10912
rect 15792 10848 15808 10912
rect 15872 10848 15888 10912
rect 15952 10848 15960 10912
rect 15640 9824 15960 10848
rect 15640 9760 15648 9824
rect 15712 9760 15728 9824
rect 15792 9760 15808 9824
rect 15872 9760 15888 9824
rect 15952 9760 15960 9824
rect 15640 8736 15960 9760
rect 15640 8672 15648 8736
rect 15712 8672 15728 8736
rect 15792 8672 15808 8736
rect 15872 8672 15888 8736
rect 15952 8672 15960 8736
rect 15640 7648 15960 8672
rect 15640 7584 15648 7648
rect 15712 7584 15728 7648
rect 15792 7584 15808 7648
rect 15872 7584 15888 7648
rect 15952 7584 15960 7648
rect 15640 6560 15960 7584
rect 15640 6496 15648 6560
rect 15712 6496 15728 6560
rect 15792 6496 15808 6560
rect 15872 6496 15888 6560
rect 15952 6496 15960 6560
rect 15640 5472 15960 6496
rect 15640 5408 15648 5472
rect 15712 5408 15728 5472
rect 15792 5408 15808 5472
rect 15872 5408 15888 5472
rect 15952 5408 15960 5472
rect 15640 4384 15960 5408
rect 15640 4320 15648 4384
rect 15712 4320 15728 4384
rect 15792 4320 15808 4384
rect 15872 4320 15888 4384
rect 15952 4320 15960 4384
rect 15640 3296 15960 4320
rect 15640 3232 15648 3296
rect 15712 3232 15728 3296
rect 15792 3232 15808 3296
rect 15872 3232 15888 3296
rect 15952 3232 15960 3296
rect 15640 2208 15960 3232
rect 15640 2144 15648 2208
rect 15712 2144 15728 2208
rect 15792 2144 15808 2208
rect 15872 2144 15888 2208
rect 15952 2144 15960 2208
rect 15640 2128 15960 2144
rect 18090 21248 18410 21808
rect 18090 21184 18098 21248
rect 18162 21184 18178 21248
rect 18242 21184 18258 21248
rect 18322 21184 18338 21248
rect 18402 21184 18410 21248
rect 18090 20160 18410 21184
rect 18090 20096 18098 20160
rect 18162 20096 18178 20160
rect 18242 20096 18258 20160
rect 18322 20096 18338 20160
rect 18402 20096 18410 20160
rect 18090 19072 18410 20096
rect 18090 19008 18098 19072
rect 18162 19008 18178 19072
rect 18242 19008 18258 19072
rect 18322 19008 18338 19072
rect 18402 19008 18410 19072
rect 18090 17984 18410 19008
rect 18090 17920 18098 17984
rect 18162 17920 18178 17984
rect 18242 17920 18258 17984
rect 18322 17920 18338 17984
rect 18402 17920 18410 17984
rect 18090 16896 18410 17920
rect 18090 16832 18098 16896
rect 18162 16832 18178 16896
rect 18242 16832 18258 16896
rect 18322 16832 18338 16896
rect 18402 16832 18410 16896
rect 18090 15808 18410 16832
rect 18090 15744 18098 15808
rect 18162 15744 18178 15808
rect 18242 15744 18258 15808
rect 18322 15744 18338 15808
rect 18402 15744 18410 15808
rect 18090 14720 18410 15744
rect 18090 14656 18098 14720
rect 18162 14656 18178 14720
rect 18242 14656 18258 14720
rect 18322 14656 18338 14720
rect 18402 14656 18410 14720
rect 18090 13632 18410 14656
rect 18090 13568 18098 13632
rect 18162 13568 18178 13632
rect 18242 13568 18258 13632
rect 18322 13568 18338 13632
rect 18402 13568 18410 13632
rect 18090 12544 18410 13568
rect 18090 12480 18098 12544
rect 18162 12480 18178 12544
rect 18242 12480 18258 12544
rect 18322 12480 18338 12544
rect 18402 12480 18410 12544
rect 18090 11456 18410 12480
rect 18090 11392 18098 11456
rect 18162 11392 18178 11456
rect 18242 11392 18258 11456
rect 18322 11392 18338 11456
rect 18402 11392 18410 11456
rect 18090 10368 18410 11392
rect 18090 10304 18098 10368
rect 18162 10304 18178 10368
rect 18242 10304 18258 10368
rect 18322 10304 18338 10368
rect 18402 10304 18410 10368
rect 18090 9280 18410 10304
rect 18090 9216 18098 9280
rect 18162 9216 18178 9280
rect 18242 9216 18258 9280
rect 18322 9216 18338 9280
rect 18402 9216 18410 9280
rect 18090 8192 18410 9216
rect 18090 8128 18098 8192
rect 18162 8128 18178 8192
rect 18242 8128 18258 8192
rect 18322 8128 18338 8192
rect 18402 8128 18410 8192
rect 18090 7104 18410 8128
rect 18090 7040 18098 7104
rect 18162 7040 18178 7104
rect 18242 7040 18258 7104
rect 18322 7040 18338 7104
rect 18402 7040 18410 7104
rect 18090 6016 18410 7040
rect 18090 5952 18098 6016
rect 18162 5952 18178 6016
rect 18242 5952 18258 6016
rect 18322 5952 18338 6016
rect 18402 5952 18410 6016
rect 18090 4928 18410 5952
rect 18090 4864 18098 4928
rect 18162 4864 18178 4928
rect 18242 4864 18258 4928
rect 18322 4864 18338 4928
rect 18402 4864 18410 4928
rect 18090 3840 18410 4864
rect 18090 3776 18098 3840
rect 18162 3776 18178 3840
rect 18242 3776 18258 3840
rect 18322 3776 18338 3840
rect 18402 3776 18410 3840
rect 18090 2752 18410 3776
rect 18090 2688 18098 2752
rect 18162 2688 18178 2752
rect 18242 2688 18258 2752
rect 18322 2688 18338 2752
rect 18402 2688 18410 2752
rect 18090 2128 18410 2688
rect 20539 21792 20859 21808
rect 20539 21728 20547 21792
rect 20611 21728 20627 21792
rect 20691 21728 20707 21792
rect 20771 21728 20787 21792
rect 20851 21728 20859 21792
rect 20539 20704 20859 21728
rect 20539 20640 20547 20704
rect 20611 20640 20627 20704
rect 20691 20640 20707 20704
rect 20771 20640 20787 20704
rect 20851 20640 20859 20704
rect 20539 19616 20859 20640
rect 20539 19552 20547 19616
rect 20611 19552 20627 19616
rect 20691 19552 20707 19616
rect 20771 19552 20787 19616
rect 20851 19552 20859 19616
rect 20539 18528 20859 19552
rect 20539 18464 20547 18528
rect 20611 18464 20627 18528
rect 20691 18464 20707 18528
rect 20771 18464 20787 18528
rect 20851 18464 20859 18528
rect 20539 17440 20859 18464
rect 20539 17376 20547 17440
rect 20611 17376 20627 17440
rect 20691 17376 20707 17440
rect 20771 17376 20787 17440
rect 20851 17376 20859 17440
rect 20539 16352 20859 17376
rect 20539 16288 20547 16352
rect 20611 16288 20627 16352
rect 20691 16288 20707 16352
rect 20771 16288 20787 16352
rect 20851 16288 20859 16352
rect 20539 15264 20859 16288
rect 20539 15200 20547 15264
rect 20611 15200 20627 15264
rect 20691 15200 20707 15264
rect 20771 15200 20787 15264
rect 20851 15200 20859 15264
rect 20539 14176 20859 15200
rect 20539 14112 20547 14176
rect 20611 14112 20627 14176
rect 20691 14112 20707 14176
rect 20771 14112 20787 14176
rect 20851 14112 20859 14176
rect 20539 13088 20859 14112
rect 20539 13024 20547 13088
rect 20611 13024 20627 13088
rect 20691 13024 20707 13088
rect 20771 13024 20787 13088
rect 20851 13024 20859 13088
rect 20539 12000 20859 13024
rect 20539 11936 20547 12000
rect 20611 11936 20627 12000
rect 20691 11936 20707 12000
rect 20771 11936 20787 12000
rect 20851 11936 20859 12000
rect 20539 10912 20859 11936
rect 20539 10848 20547 10912
rect 20611 10848 20627 10912
rect 20691 10848 20707 10912
rect 20771 10848 20787 10912
rect 20851 10848 20859 10912
rect 20539 9824 20859 10848
rect 20539 9760 20547 9824
rect 20611 9760 20627 9824
rect 20691 9760 20707 9824
rect 20771 9760 20787 9824
rect 20851 9760 20859 9824
rect 20539 8736 20859 9760
rect 20539 8672 20547 8736
rect 20611 8672 20627 8736
rect 20691 8672 20707 8736
rect 20771 8672 20787 8736
rect 20851 8672 20859 8736
rect 20539 7648 20859 8672
rect 20539 7584 20547 7648
rect 20611 7584 20627 7648
rect 20691 7584 20707 7648
rect 20771 7584 20787 7648
rect 20851 7584 20859 7648
rect 20539 6560 20859 7584
rect 20539 6496 20547 6560
rect 20611 6496 20627 6560
rect 20691 6496 20707 6560
rect 20771 6496 20787 6560
rect 20851 6496 20859 6560
rect 20539 5472 20859 6496
rect 20539 5408 20547 5472
rect 20611 5408 20627 5472
rect 20691 5408 20707 5472
rect 20771 5408 20787 5472
rect 20851 5408 20859 5472
rect 20539 4384 20859 5408
rect 20539 4320 20547 4384
rect 20611 4320 20627 4384
rect 20691 4320 20707 4384
rect 20771 4320 20787 4384
rect 20851 4320 20859 4384
rect 20539 3296 20859 4320
rect 21219 3500 21285 3501
rect 21219 3436 21220 3500
rect 21284 3436 21285 3500
rect 21219 3435 21285 3436
rect 20539 3232 20547 3296
rect 20611 3232 20627 3296
rect 20691 3232 20707 3296
rect 20771 3232 20787 3296
rect 20851 3232 20859 3296
rect 20539 2208 20859 3232
rect 21222 3229 21282 3435
rect 21219 3228 21285 3229
rect 21219 3164 21220 3228
rect 21284 3164 21285 3228
rect 21219 3163 21285 3164
rect 20539 2144 20547 2208
rect 20611 2144 20627 2208
rect 20691 2144 20707 2208
rect 20771 2144 20787 2208
rect 20851 2144 20859 2208
rect 20539 2128 20859 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1662439860
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1662439860
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1662439860
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1662439860
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1662439860
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105
timestamp 1662439860
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1662439860
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1662439860
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1662439860
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1662439860
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1662439860
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155
timestamp 1662439860
transform 1 0 15364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1662439860
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1662439860
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1662439860
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_183 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 17940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1662439860
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1662439860
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1662439860
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_203
timestamp 1662439860
transform 1 0 19780 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_209
timestamp 1662439860
transform 1 0 20332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1662439860
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1662439860
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1662439860
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_42
timestamp 1662439860
transform 1 0 4968 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1662439860
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1662439860
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_79
timestamp 1662439860
transform 1 0 8372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1662439860
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1662439860
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1662439860
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1662439860
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1662439860
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1662439860
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1662439860
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1662439860
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1662439860
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1662439860
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1662439860
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1662439860
transform 1 0 20240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1662439860
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1662439860
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_17
timestamp 1662439860
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1662439860
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1662439860
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1662439860
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_63
timestamp 1662439860
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1662439860
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1662439860
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1662439860
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_97
timestamp 1662439860
transform 1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_124
timestamp 1662439860
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1662439860
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1662439860
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp 1662439860
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1662439860
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1662439860
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1662439860
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1662439860
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_203
timestamp 1662439860
transform 1 0 19780 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1662439860
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1662439860
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_28
timestamp 1662439860
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1662439860
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1662439860
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1662439860
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_62
timestamp 1662439860
transform 1 0 6808 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_74
timestamp 1662439860
transform 1 0 7912 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_96
timestamp 1662439860
transform 1 0 9936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1662439860
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1662439860
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1662439860
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1662439860
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1662439860
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1662439860
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1662439860
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1662439860
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_201
timestamp 1662439860
transform 1 0 19596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_209
timestamp 1662439860
transform 1 0 20332 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1662439860
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1662439860
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1662439860
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_37
timestamp 1662439860
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_43
timestamp 1662439860
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_55
timestamp 1662439860
transform 1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1662439860
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1662439860
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1662439860
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_92
timestamp 1662439860
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_99
timestamp 1662439860
transform 1 0 10212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_111
timestamp 1662439860
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_123
timestamp 1662439860
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1662439860
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1662439860
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp 1662439860
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_149
timestamp 1662439860
transform 1 0 14812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1662439860
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_178
timestamp 1662439860
transform 1 0 17480 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1662439860
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1662439860
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1662439860
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1662439860
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1662439860
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1662439860
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1662439860
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1662439860
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1662439860
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1662439860
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_64
timestamp 1662439860
transform 1 0 6992 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp 1662439860
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1662439860
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_100
timestamp 1662439860
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1662439860
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1662439860
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 1662439860
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1662439860
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1662439860
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_195
timestamp 1662439860
transform 1 0 19044 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_203
timestamp 1662439860
transform 1 0 19780 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1662439860
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1662439860
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1662439860
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1662439860
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1662439860
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1662439860
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_60
timestamp 1662439860
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1662439860
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1662439860
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1662439860
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1662439860
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_95
timestamp 1662439860
transform 1 0 9844 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1662439860
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1662439860
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1662439860
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp 1662439860
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1662439860
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_167
timestamp 1662439860
transform 1 0 16468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1662439860
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1662439860
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1662439860
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_209
timestamp 1662439860
transform 1 0 20332 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1662439860
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1662439860
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1662439860
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_22
timestamp 1662439860
transform 1 0 3128 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1662439860
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_42
timestamp 1662439860
transform 1 0 4968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1662439860
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1662439860
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1662439860
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_74
timestamp 1662439860
transform 1 0 7912 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1662439860
transform 1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1662439860
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_99
timestamp 1662439860
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1662439860
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1662439860
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1662439860
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_142
timestamp 1662439860
transform 1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1662439860
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1662439860
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_191
timestamp 1662439860
transform 1 0 18676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_203
timestamp 1662439860
transform 1 0 19780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_209
timestamp 1662439860
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1662439860
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1662439860
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1662439860
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1662439860
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1662439860
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_34
timestamp 1662439860
transform 1 0 4232 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_69
timestamp 1662439860
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1662439860
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1662439860
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_90
timestamp 1662439860
transform 1 0 9384 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_94
timestamp 1662439860
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_98
timestamp 1662439860
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_113
timestamp 1662439860
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_125
timestamp 1662439860
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1662439860
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1662439860
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1662439860
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_157
timestamp 1662439860
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_161
timestamp 1662439860
transform 1 0 15916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_173
timestamp 1662439860
transform 1 0 17020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp 1662439860
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1662439860
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1662439860
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1662439860
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1662439860
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1662439860
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_25
timestamp 1662439860
transform 1 0 3404 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 1662439860
transform 1 0 4140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_40
timestamp 1662439860
transform 1 0 4784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1662439860
transform 1 0 5520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1662439860
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1662439860
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp 1662439860
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1662439860
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_84
timestamp 1662439860
transform 1 0 8832 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1662439860
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1662439860
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_118
timestamp 1662439860
transform 1 0 11960 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_130
timestamp 1662439860
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_142
timestamp 1662439860
transform 1 0 14168 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_148
timestamp 1662439860
transform 1 0 14720 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_152
timestamp 1662439860
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1662439860
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1662439860
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1662439860
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1662439860
transform 1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1662439860
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1662439860
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1662439860
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1662439860
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1662439860
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_47
timestamp 1662439860
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_59
timestamp 1662439860
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1662439860
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1662439860
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp 1662439860
transform 1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1662439860
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_131
timestamp 1662439860
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1662439860
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1662439860
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1662439860
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1662439860
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1662439860
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_181
timestamp 1662439860
transform 1 0 17756 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1662439860
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1662439860
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1662439860
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1662439860
transform 1 0 19688 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1662439860
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_20
timestamp 1662439860
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_28
timestamp 1662439860
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1662439860
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1662439860
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1662439860
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_63
timestamp 1662439860
transform 1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_72
timestamp 1662439860
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_96
timestamp 1662439860
transform 1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1662439860
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1662439860
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1662439860
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1662439860
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1662439860
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1662439860
transform 1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1662439860
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1662439860
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1662439860
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1662439860
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_198
timestamp 1662439860
transform 1 0 19320 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1662439860
transform 1 0 20240 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1662439860
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_15
timestamp 1662439860
transform 1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1662439860
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1662439860
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1662439860
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1662439860
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_42
timestamp 1662439860
transform 1 0 4968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1662439860
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1662439860
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1662439860
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1662439860
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1662439860
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_96
timestamp 1662439860
transform 1 0 9936 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_108
timestamp 1662439860
transform 1 0 11040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1662439860
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1662439860
transform 1 0 12880 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1662439860
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1662439860
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1662439860
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_149
timestamp 1662439860
transform 1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_172
timestamp 1662439860
transform 1 0 16928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_179
timestamp 1662439860
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_183
timestamp 1662439860
transform 1 0 17940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1662439860
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1662439860
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1662439860
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_203
timestamp 1662439860
transform 1 0 19780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_209
timestamp 1662439860
transform 1 0 20332 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1662439860
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_13
timestamp 1662439860
transform 1 0 2300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1662439860
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_41
timestamp 1662439860
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1662439860
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1662439860
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_65
timestamp 1662439860
transform 1 0 7084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_77
timestamp 1662439860
transform 1 0 8188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1662439860
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1662439860
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1662439860
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1662439860
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1662439860
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1662439860
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1662439860
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1662439860
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1662439860
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1662439860
transform 1 0 18032 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1662439860
transform 1 0 20240 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1662439860
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1662439860
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1662439860
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1662439860
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1662439860
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1662439860
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_65
timestamp 1662439860
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_73
timestamp 1662439860
transform 1 0 7820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1662439860
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1662439860
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1662439860
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1662439860
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_104
timestamp 1662439860
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1662439860
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_122
timestamp 1662439860
transform 1 0 12328 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1662439860
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1662439860
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_163
timestamp 1662439860
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1662439860
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1662439860
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1662439860
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1662439860
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 1662439860
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_208
timestamp 1662439860
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1662439860
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_8
timestamp 1662439860
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1662439860
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1662439860
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1662439860
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1662439860
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_69
timestamp 1662439860
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1662439860
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1662439860
transform 1 0 10396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1662439860
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1662439860
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1662439860
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1662439860
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1662439860
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1662439860
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1662439860
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1662439860
transform 1 0 20240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1662439860
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_8
timestamp 1662439860
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1662439860
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1662439860
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_39
timestamp 1662439860
transform 1 0 4692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_48
timestamp 1662439860
transform 1 0 5520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_54
timestamp 1662439860
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1662439860
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1662439860
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1662439860
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1662439860
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1662439860
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1662439860
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_114
timestamp 1662439860
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_126
timestamp 1662439860
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1662439860
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1662439860
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1662439860
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_159
timestamp 1662439860
transform 1 0 15732 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_176
timestamp 1662439860
transform 1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_183
timestamp 1662439860
transform 1 0 17940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1662439860
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1662439860
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1662439860
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1662439860
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1662439860
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_23
timestamp 1662439860
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1662439860
transform 1 0 3772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_41
timestamp 1662439860
transform 1 0 4876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1662439860
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1662439860
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1662439860
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_63
timestamp 1662439860
transform 1 0 6900 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_75
timestamp 1662439860
transform 1 0 8004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_87
timestamp 1662439860
transform 1 0 9108 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1662439860
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1662439860
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1662439860
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_119
timestamp 1662439860
transform 1 0 12052 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1662439860
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1662439860
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1662439860
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1662439860
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1662439860
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_188
timestamp 1662439860
transform 1 0 18400 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_200
timestamp 1662439860
transform 1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1662439860
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1662439860
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_8
timestamp 1662439860
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1662439860
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1662439860
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1662439860
transform 1 0 4784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1662439860
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1662439860
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_61
timestamp 1662439860
transform 1 0 6716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_67
timestamp 1662439860
transform 1 0 7268 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_71
timestamp 1662439860
transform 1 0 7636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1662439860
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1662439860
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_107
timestamp 1662439860
transform 1 0 10948 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1662439860
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1662439860
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1662439860
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1662439860
transform 1 0 14628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_173
timestamp 1662439860
transform 1 0 17020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1662439860
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1662439860
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1662439860
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1662439860
transform 1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1662439860
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1662439860
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_19
timestamp 1662439860
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1662439860
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1662439860
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1662439860
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1662439860
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1662439860
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_86
timestamp 1662439860
transform 1 0 9016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1662439860
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1662439860
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1662439860
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_120
timestamp 1662439860
transform 1 0 12144 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1662439860
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_138
timestamp 1662439860
transform 1 0 13800 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1662439860
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1662439860
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1662439860
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_181
timestamp 1662439860
transform 1 0 17756 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_187
timestamp 1662439860
transform 1 0 18308 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1662439860
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1662439860
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_12
timestamp 1662439860
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1662439860
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1662439860
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_41
timestamp 1662439860
transform 1 0 4876 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_47
timestamp 1662439860
transform 1 0 5428 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_68
timestamp 1662439860
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1662439860
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1662439860
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1662439860
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_103
timestamp 1662439860
transform 1 0 10580 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1662439860
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1662439860
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_128
timestamp 1662439860
transform 1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1662439860
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1662439860
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1662439860
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1662439860
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1662439860
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1662439860
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1662439860
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1662439860
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp 1662439860
transform 1 0 20240 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1662439860
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_8
timestamp 1662439860
transform 1 0 1840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1662439860
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_40
timestamp 1662439860
transform 1 0 4784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1662439860
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1662439860
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1662439860
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_65
timestamp 1662439860
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_69
timestamp 1662439860
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_84
timestamp 1662439860
transform 1 0 8832 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1662439860
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1662439860
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_118
timestamp 1662439860
transform 1 0 11960 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_144
timestamp 1662439860
transform 1 0 14352 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_156
timestamp 1662439860
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1662439860
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_181
timestamp 1662439860
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_187
timestamp 1662439860
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_208
timestamp 1662439860
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1662439860
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_9
timestamp 1662439860
transform 1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1662439860
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1662439860
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1662439860
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1662439860
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1662439860
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_66
timestamp 1662439860
transform 1 0 7176 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1662439860
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1662439860
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1662439860
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1662439860
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_116
timestamp 1662439860
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1662439860
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1662439860
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1662439860
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_163
timestamp 1662439860
transform 1 0 16100 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1662439860
transform 1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1662439860
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1662439860
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1662439860
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 1662439860
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1662439860
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_8
timestamp 1662439860
transform 1 0 1840 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_20
timestamp 1662439860
transform 1 0 2944 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_32
timestamp 1662439860
transform 1 0 4048 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_44
timestamp 1662439860
transform 1 0 5152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1662439860
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1662439860
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1662439860
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_65
timestamp 1662439860
transform 1 0 7084 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_73
timestamp 1662439860
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_85
timestamp 1662439860
transform 1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1662439860
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1662439860
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1662439860
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1662439860
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1662439860
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_121
timestamp 1662439860
transform 1 0 12236 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_133
timestamp 1662439860
transform 1 0 13340 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_139
timestamp 1662439860
transform 1 0 13892 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_143
timestamp 1662439860
transform 1 0 14260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_155
timestamp 1662439860
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1662439860
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1662439860
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_181
timestamp 1662439860
transform 1 0 17756 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_187
timestamp 1662439860
transform 1 0 18308 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_208
timestamp 1662439860
transform 1 0 20240 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1662439860
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1662439860
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_11
timestamp 1662439860
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1662439860
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1662439860
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1662439860
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1662439860
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1662439860
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1662439860
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_72
timestamp 1662439860
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1662439860
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1662439860
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1662439860
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_102
timestamp 1662439860
transform 1 0 10488 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_123
timestamp 1662439860
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1662439860
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1662439860
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1662439860
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_149
timestamp 1662439860
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1662439860
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1662439860
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1662439860
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1662439860
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_208
timestamp 1662439860
transform 1 0 20240 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1662439860
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_26
timestamp 1662439860
transform 1 0 3496 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_38
timestamp 1662439860
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1662439860
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1662439860
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1662439860
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_67
timestamp 1662439860
transform 1 0 7268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_74
timestamp 1662439860
transform 1 0 7912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_78
timestamp 1662439860
transform 1 0 8280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1662439860
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1662439860
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1662439860
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1662439860
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1662439860
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_130
timestamp 1662439860
transform 1 0 13064 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_138
timestamp 1662439860
transform 1 0 13800 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_147
timestamp 1662439860
transform 1 0 14628 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1662439860
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1662439860
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1662439860
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1662439860
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_175
timestamp 1662439860
transform 1 0 17204 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp 1662439860
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_208
timestamp 1662439860
transform 1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1662439860
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_16
timestamp 1662439860
transform 1 0 2576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1662439860
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1662439860
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1662439860
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_36
timestamp 1662439860
transform 1 0 4416 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_43
timestamp 1662439860
transform 1 0 5060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_55
timestamp 1662439860
transform 1 0 6164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1662439860
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1662439860
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1662439860
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1662439860
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_124
timestamp 1662439860
transform 1 0 12512 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_130
timestamp 1662439860
transform 1 0 13064 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1662439860
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1662439860
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1662439860
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1662439860
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1662439860
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1662439860
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1662439860
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1662439860
transform 1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1662439860
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_25
timestamp 1662439860
transform 1 0 3404 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_32
timestamp 1662439860
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1662439860
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1662439860
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_68
timestamp 1662439860
transform 1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_75
timestamp 1662439860
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_87
timestamp 1662439860
transform 1 0 9108 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_94
timestamp 1662439860
transform 1 0 9752 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1662439860
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1662439860
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_121
timestamp 1662439860
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_127
timestamp 1662439860
transform 1 0 12788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_139
timestamp 1662439860
transform 1 0 13892 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1662439860
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1662439860
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1662439860
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_174
timestamp 1662439860
transform 1 0 17112 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_202
timestamp 1662439860
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1662439860
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_17
timestamp 1662439860
transform 1 0 2668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1662439860
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1662439860
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1662439860
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_63
timestamp 1662439860
transform 1 0 6900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_67
timestamp 1662439860
transform 1 0 7268 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_71
timestamp 1662439860
transform 1 0 7636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1662439860
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1662439860
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_94
timestamp 1662439860
transform 1 0 9752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_100
timestamp 1662439860
transform 1 0 10304 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_105
timestamp 1662439860
transform 1 0 10764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_113
timestamp 1662439860
transform 1 0 11500 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1662439860
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1662439860
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_150
timestamp 1662439860
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_162
timestamp 1662439860
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1662439860
transform 1 0 16744 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_175
timestamp 1662439860
transform 1 0 17204 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_184
timestamp 1662439860
transform 1 0 18032 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1662439860
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1662439860
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1662439860
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_208
timestamp 1662439860
transform 1 0 20240 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1662439860
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1662439860
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_16
timestamp 1662439860
transform 1 0 2576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1662439860
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1662439860
transform 1 0 4048 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1662439860
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1662439860
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_79
timestamp 1662439860
transform 1 0 8372 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_87
timestamp 1662439860
transform 1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1662439860
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1662439860
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_119
timestamp 1662439860
transform 1 0 12052 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_126
timestamp 1662439860
transform 1 0 12696 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_138
timestamp 1662439860
transform 1 0 13800 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_144
timestamp 1662439860
transform 1 0 14352 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1662439860
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1662439860
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_176
timestamp 1662439860
transform 1 0 17296 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_202
timestamp 1662439860
transform 1 0 19688 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1662439860
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1662439860
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1662439860
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1662439860
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1662439860
transform 1 0 5796 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_59
timestamp 1662439860
transform 1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1662439860
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1662439860
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1662439860
transform 1 0 10028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1662439860
transform 1 0 10580 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_125
timestamp 1662439860
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1662439860
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1662439860
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_153
timestamp 1662439860
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1662439860
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1662439860
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1662439860
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1662439860
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1662439860
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_203
timestamp 1662439860
transform 1 0 19780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_208
timestamp 1662439860
transform 1 0 20240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1662439860
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1662439860
transform 1 0 2116 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1662439860
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1662439860
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1662439860
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1662439860
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_63
timestamp 1662439860
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_84
timestamp 1662439860
transform 1 0 8832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1662439860
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1662439860
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1662439860
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1662439860
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1662439860
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1662439860
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1662439860
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1662439860
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1662439860
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1662439860
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_185
timestamp 1662439860
transform 1 0 18124 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1662439860
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1662439860
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_15
timestamp 1662439860
transform 1 0 2484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1662439860
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1662439860
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1662439860
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1662439860
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1662439860
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1662439860
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1662439860
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp 1662439860
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_105
timestamp 1662439860
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_128
timestamp 1662439860
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1662439860
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1662439860
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1662439860
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1662439860
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1662439860
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_204
timestamp 1662439860
transform 1 0 19872 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1662439860
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_9
timestamp 1662439860
transform 1 0 1932 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1662439860
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_19
timestamp 1662439860
transform 1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_43
timestamp 1662439860
transform 1 0 5060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1662439860
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1662439860
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_63
timestamp 1662439860
transform 1 0 6900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_70
timestamp 1662439860
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_95
timestamp 1662439860
transform 1 0 9844 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1662439860
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1662439860
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1662439860
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1662439860
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1662439860
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1662439860
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1662439860
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1662439860
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_200
timestamp 1662439860
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_208
timestamp 1662439860
transform 1 0 20240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1662439860
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_9
timestamp 1662439860
transform 1 0 1932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_15
timestamp 1662439860
transform 1 0 2484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1662439860
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1662439860
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_37
timestamp 1662439860
transform 1 0 4508 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_60
timestamp 1662439860
transform 1 0 6624 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_68
timestamp 1662439860
transform 1 0 7360 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1662439860
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1662439860
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1662439860
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_97
timestamp 1662439860
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_118
timestamp 1662439860
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_126
timestamp 1662439860
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1662439860
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1662439860
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_153
timestamp 1662439860
transform 1 0 15180 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1662439860
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_183
timestamp 1662439860
transform 1 0 17940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1662439860
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1662439860
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1662439860
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_208
timestamp 1662439860
transform 1 0 20240 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1662439860
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_13
timestamp 1662439860
transform 1 0 2300 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_21
timestamp 1662439860
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_26
timestamp 1662439860
transform 1 0 3496 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_29
timestamp 1662439860
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_41
timestamp 1662439860
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1662439860
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1662439860
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1662439860
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_69
timestamp 1662439860
transform 1 0 7452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_77
timestamp 1662439860
transform 1 0 8188 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_82
timestamp 1662439860
transform 1 0 8648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_85
timestamp 1662439860
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_97
timestamp 1662439860
transform 1 0 10028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_105
timestamp 1662439860
transform 1 0 10764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1662439860
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1662439860
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1662439860
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_137
timestamp 1662439860
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_141
timestamp 1662439860
transform 1 0 14076 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1662439860
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_155
timestamp 1662439860
transform 1 0 15364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 1662439860
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1662439860
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_175
timestamp 1662439860
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_183
timestamp 1662439860
transform 1 0 17940 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1662439860
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1662439860
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1662439860
transform 1 0 19228 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_203
timestamp 1662439860
transform 1 0 19780 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_209
timestamp 1662439860
transform 1 0 20332 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1662439860
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1662439860
transform -1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1662439860
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1662439860
transform -1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1662439860
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1662439860
transform -1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1662439860
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1662439860
transform -1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1662439860
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1662439860
transform -1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1662439860
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1662439860
transform -1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1662439860
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1662439860
transform -1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1662439860
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1662439860
transform -1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1662439860
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1662439860
transform -1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1662439860
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1662439860
transform -1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1662439860
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1662439860
transform -1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1662439860
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1662439860
transform -1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1662439860
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1662439860
transform -1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1662439860
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1662439860
transform -1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1662439860
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1662439860
transform -1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1662439860
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1662439860
transform -1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1662439860
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1662439860
transform -1 0 20700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1662439860
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1662439860
transform -1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1662439860
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1662439860
transform -1 0 20700 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1662439860
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1662439860
transform -1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1662439860
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1662439860
transform -1 0 20700 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1662439860
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1662439860
transform -1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1662439860
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1662439860
transform -1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1662439860
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1662439860
transform -1 0 20700 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1662439860
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1662439860
transform -1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1662439860
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1662439860
transform -1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1662439860
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1662439860
transform -1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1662439860
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1662439860
transform -1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1662439860
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1662439860
transform -1 0 20700 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1662439860
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1662439860
transform -1 0 20700 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1662439860
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1662439860
transform -1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1662439860
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1662439860
transform -1 0 20700 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1662439860
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1662439860
transform -1 0 20700 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1662439860
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1662439860
transform -1 0 20700 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1662439860
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1662439860
transform -1 0 20700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1662439860
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1662439860
transform -1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1662439860
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1662439860
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1662439860
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1662439860
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1662439860
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1662439860
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1662439860
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1662439860
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1662439860
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1662439860
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1662439860
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1662439860
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1662439860
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1662439860
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1662439860
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1662439860
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1662439860
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1662439860
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1662439860
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1662439860
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1662439860
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1662439860
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1662439860
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1662439860
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1662439860
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1662439860
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1662439860
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1662439860
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1662439860
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1662439860
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1662439860
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1662439860
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1662439860
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1662439860
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1662439860
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1662439860
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1662439860
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1662439860
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1662439860
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1662439860
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1662439860
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1662439860
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1662439860
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1662439860
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1662439860
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1662439860
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1662439860
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1662439860
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1662439860
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1662439860
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1662439860
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1662439860
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1662439860
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1662439860
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1662439860
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1662439860
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1662439860
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1662439860
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1662439860
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1662439860
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1662439860
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1662439860
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1662439860
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1662439860
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1662439860
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1662439860
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1662439860
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1662439860
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1662439860
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1662439860
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1662439860
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1662439860
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1662439860
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1662439860
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1662439860
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1662439860
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1662439860
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1662439860
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1662439860
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1662439860
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1662439860
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1662439860
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1662439860
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1662439860
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1662439860
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1662439860
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1662439860
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1662439860
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1662439860
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1662439860
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1662439860
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1662439860
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1662439860
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1662439860
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1662439860
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1662439860
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1662439860
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1662439860
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1662439860
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1662439860
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1662439860
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1662439860
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1662439860
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1662439860
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1662439860
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1662439860
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1662439860
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1662439860
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1662439860
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1662439860
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1662439860
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1662439860
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1662439860
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1662439860
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1662439860
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1662439860
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1662439860
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1662439860
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1662439860
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1662439860
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1662439860
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1662439860
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1662439860
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1662439860
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1662439860
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1662439860
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1662439860
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1662439860
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1662439860
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1662439860
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1662439860
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1662439860
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  fanout52 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9384 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 11132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 1662439860
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1662439860
transform 1 0 14904 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1662439860
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1662439860
transform -1 0 16376 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout58 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 17756 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1662439860
transform -1 0 19780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 1662439860
transform -1 0 7084 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout61 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1662439860
transform -1 0 6072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 1662439860
transform -1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 1662439860
transform -1 0 14628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 1662439860
transform -1 0 12052 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1662439860
transform 1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout67
timestamp 1662439860
transform -1 0 2944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 1662439860
transform -1 0 2944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1662439860
transform -1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1662439860
transform -1 0 20240 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 1662439860
transform -1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 1662439860
transform 1 0 18584 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp 1662439860
transform -1 0 7360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout74
timestamp 1662439860
transform -1 0 13800 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1662439860
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1662439860
transform -1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1662439860
transform -1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1662439860
transform -1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1662439860
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1662439860
transform -1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1662439860
transform -1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1662439860
transform -1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1662439860
transform -1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1662439860
transform -1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1662439860
transform -1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1662439860
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1662439860
transform 1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1662439860
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1662439860
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1662439860
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1662439860
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1662439860
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1662439860
transform -1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1662439860
transform -1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1662439860
transform -1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1662439860
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1662439860
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1662439860
transform -1 0 18952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1662439860
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1662439860
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1662439860
transform -1 0 15364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1662439860
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1662439860
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1662439860
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1662439860
transform -1 0 6072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1662439860
transform -1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1662439860
transform 1 0 19412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1662439860
transform 1 0 17572 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1662439860
transform -1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1662439860
transform -1 0 11224 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1662439860
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1662439860
transform -1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1662439860
transform -1 0 3496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1662439860
transform -1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1662439860
transform -1 0 18952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1662439860
transform 1 0 19872 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1662439860
transform 1 0 16836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1662439860
transform 1 0 14996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1662439860
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1662439860
transform 1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1662439860
transform 1 0 7084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1662439860
transform 1 0 5704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1662439860
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1662439860
transform -1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  x1_x1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 10028 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x2
timestamp 1662439860
transform 1 0 10580 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x3
timestamp 1662439860
transform 1 0 5336 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x4
timestamp 1662439860
transform 1 0 5520 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x5
timestamp 1662439860
transform 1 0 6532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x6
timestamp 1662439860
transform 1 0 6164 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x7
timestamp 1662439860
transform 1 0 6808 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x8
timestamp 1662439860
transform 1 0 8096 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x9
timestamp 1662439860
transform 1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x10
timestamp 1662439860
transform 1 0 10672 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x11
timestamp 1662439860
transform 1 0 12512 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x12
timestamp 1662439860
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x13
timestamp 1662439860
transform 1 0 15088 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x14
timestamp 1662439860
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  x1_x15
timestamp 1662439860
transform -1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x16
timestamp 1662439860
transform -1 0 7268 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x17
timestamp 1662439860
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x18
timestamp 1662439860
transform -1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x19
timestamp 1662439860
transform 1 0 10580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x20
timestamp 1662439860
transform -1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x21
timestamp 1662439860
transform 1 0 5520 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x22
timestamp 1662439860
transform 1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x23
timestamp 1662439860
transform -1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x24
timestamp 1662439860
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x25
timestamp 1662439860
transform -1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x26
timestamp 1662439860
transform -1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x27
timestamp 1662439860
transform -1 0 6900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  x1_x28
timestamp 1662439860
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x29
timestamp 1662439860
transform -1 0 10120 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x30
timestamp 1662439860
transform -1 0 4968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x1_x31
timestamp 1662439860
transform 1 0 6808 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x1_x32
timestamp 1662439860
transform 1 0 8372 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  x1_x33
timestamp 1662439860
transform -1 0 5612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x1_x34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3772 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x1_x35 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3956 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  x1_x36_75 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 7636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x1_x36 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x37
timestamp 1662439860
transform -1 0 5060 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x38
timestamp 1662439860
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x39
timestamp 1662439860
transform -1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x40
timestamp 1662439860
transform -1 0 13064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x41
timestamp 1662439860
transform 1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x42
timestamp 1662439860
transform -1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x43
timestamp 1662439860
transform -1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x44
timestamp 1662439860
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x45
timestamp 1662439860
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x46
timestamp 1662439860
transform -1 0 8004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x47
timestamp 1662439860
transform -1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x48
timestamp 1662439860
transform -1 0 6072 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x49
timestamp 1662439860
transform -1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x50
timestamp 1662439860
transform -1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x51
timestamp 1662439860
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x52
timestamp 1662439860
transform -1 0 7728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x53
timestamp 1662439860
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x54
timestamp 1662439860
transform -1 0 10580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x55
timestamp 1662439860
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x56
timestamp 1662439860
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x57
timestamp 1662439860
transform 1 0 15364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x58
timestamp 1662439860
transform -1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  x1_x59
timestamp 1662439860
transform -1 0 6900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x60
timestamp 1662439860
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x61
timestamp 1662439860
transform -1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x62
timestamp 1662439860
transform -1 0 12512 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x63
timestamp 1662439860
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x64
timestamp 1662439860
transform -1 0 12144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x65
timestamp 1662439860
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x66
timestamp 1662439860
transform -1 0 12420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x67
timestamp 1662439860
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x68
timestamp 1662439860
transform 1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  x1_x69
timestamp 1662439860
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  x1_x70
timestamp 1662439860
transform -1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x71
timestamp 1662439860
transform -1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x72
timestamp 1662439860
transform -1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x73
timestamp 1662439860
transform -1 0 17572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x74
timestamp 1662439860
transform -1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x75
timestamp 1662439860
transform -1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x76
timestamp 1662439860
transform -1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x77
timestamp 1662439860
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x1_x78
timestamp 1662439860
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x2
timestamp 1662439860
transform -1 0 18492 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__fa_1  x3_x62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 17296 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x3_x64
timestamp 1662439860
transform 1 0 17020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x3_x65
timestamp 1662439860
transform 1 0 17388 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  x3_x67
timestamp 1662439860
transform 1 0 18400 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x3_x68
timestamp 1662439860
transform 1 0 18400 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__fa_1  x3_x69
timestamp 1662439860
transform 1 0 16928 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  x3_x70
timestamp 1662439860
transform 1 0 18400 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x3_x71
timestamp 1662439860
transform 1 0 18400 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__fa_1  x3_x72
timestamp 1662439860
transform 1 0 15824 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x3_x73
timestamp 1662439860
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  x3_x74
timestamp 1662439860
transform 1 0 18400 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x3_x75
timestamp 1662439860
transform 1 0 18400 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fa_1  x3_x76
timestamp 1662439860
transform 1 0 14996 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  x3_x77
timestamp 1662439860
transform 1 0 14904 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  x3_x78
timestamp 1662439860
transform 1 0 17204 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x3_x79
timestamp 1662439860
transform 1 0 17756 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x3_x80
timestamp 1662439860
transform 1 0 18400 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x3_x81
timestamp 1662439860
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x3_x82
timestamp 1662439860
transform 1 0 16928 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x1
timestamp 1662439860
transform 1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x2
timestamp 1662439860
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  x4_x3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 11684 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  x4_x4
timestamp 1662439860
transform 1 0 16468 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x5
timestamp 1662439860
transform 1 0 15088 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  x4_x6
timestamp 1662439860
transform 1 0 13616 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  x4_x7
timestamp 1662439860
transform 1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x8
timestamp 1662439860
transform 1 0 15180 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x9
timestamp 1662439860
transform 1 0 14260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  x4_x10
timestamp 1662439860
transform 1 0 5336 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  x4_x11
timestamp 1662439860
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x12
timestamp 1662439860
transform 1 0 11684 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x13
timestamp 1662439860
transform 1 0 12328 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x14
timestamp 1662439860
transform 1 0 13892 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x15
timestamp 1662439860
transform 1 0 16836 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__and2_0  x4_x16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 13156 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x17
timestamp 1662439860
transform 1 0 11868 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x18
timestamp 1662439860
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x19
timestamp 1662439860
transform -1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x20
timestamp 1662439860
transform 1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x21 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x4_x22
timestamp 1662439860
transform 1 0 16836 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_0  x4_x23
timestamp 1662439860
transform 1 0 17572 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x24_x1
timestamp 1662439860
transform -1 0 17296 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x24_x2
timestamp 1662439860
transform 1 0 17480 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x24_x3
timestamp 1662439860
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x25
timestamp 1662439860
transform 1 0 17848 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__and2_0  x4_x26
timestamp 1662439860
transform 1 0 12420 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  x4_x27
timestamp 1662439860
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  x4_x28
timestamp 1662439860
transform 1 0 15456 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__xor2_1  x4_x29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14260 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  x4_x30_x1
timestamp 1662439860
transform -1 0 15732 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x30_x2
timestamp 1662439860
transform 1 0 15732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x30_x3
timestamp 1662439860
transform -1 0 16376 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  x4_x31
timestamp 1662439860
transform 1 0 13156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  x4_x32
timestamp 1662439860
transform 1 0 10580 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_0  x4_x33
timestamp 1662439860
transform -1 0 9568 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x34_x1
timestamp 1662439860
transform 1 0 11316 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x34_x2
timestamp 1662439860
transform 1 0 10672 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x34_x3
timestamp 1662439860
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x35
timestamp 1662439860
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__and2_0  x4_x36
timestamp 1662439860
transform 1 0 6532 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  x4_x37
timestamp 1662439860
transform 1 0 8188 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  x4_x38
timestamp 1662439860
transform 1 0 9292 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_0  x4_x39_x1
timestamp 1662439860
transform 1 0 10396 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x39_x2
timestamp 1662439860
transform 1 0 11684 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x39_x3
timestamp 1662439860
transform 1 0 9844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  x4_x40
timestamp 1662439860
transform 1 0 8004 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  x4_x41
timestamp 1662439860
transform 1 0 13892 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x4_x42
timestamp 1662439860
transform 1 0 7268 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  x4_x43
timestamp 1662439860
transform 1 0 8004 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  x4_x44_x1
timestamp 1662439860
transform -1 0 10856 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x44_x2
timestamp 1662439860
transform 1 0 11040 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x44_x3
timestamp 1662439860
transform 1 0 9292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  x4_x45
timestamp 1662439860
transform 1 0 7544 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  x4_x46
timestamp 1662439860
transform 1 0 19412 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x47
timestamp 1662439860
transform 1 0 4324 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  x4_x48
timestamp 1662439860
transform 1 0 14444 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 16376 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x50 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 15272 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x51
timestamp 1662439860
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x52
timestamp 1662439860
transform 1 0 14628 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x53
timestamp 1662439860
transform 1 0 13892 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x54
timestamp 1662439860
transform 1 0 9108 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x55
timestamp 1662439860
transform 1 0 9936 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x56
timestamp 1662439860
transform 1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x57
timestamp 1662439860
transform 1 0 9108 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x58
timestamp 1662439860
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x59
timestamp 1662439860
transform 1 0 9936 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x60
timestamp 1662439860
transform 1 0 8556 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x61
timestamp 1662439860
transform 1 0 1564 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  x4_x62
timestamp 1662439860
transform 1 0 2852 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x63
timestamp 1662439860
transform 1 0 9936 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  x4_x64
timestamp 1662439860
transform -1 0 2484 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  x4_x65
timestamp 1662439860
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x66
timestamp 1662439860
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x67
timestamp 1662439860
transform 1 0 6532 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x68
timestamp 1662439860
transform 1 0 6348 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x69
timestamp 1662439860
transform 1 0 5060 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x70
timestamp 1662439860
transform 1 0 5060 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x71
timestamp 1662439860
transform 1 0 4048 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x72
timestamp 1662439860
transform 1 0 3956 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x73
timestamp 1662439860
transform -1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x74
timestamp 1662439860
transform 1 0 2944 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x4_x75
timestamp 1662439860
transform 1 0 3036 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x76
timestamp 1662439860
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x77
timestamp 1662439860
transform -1 0 3680 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x4_x78
timestamp 1662439860
transform 1 0 2208 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x79
timestamp 1662439860
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x80
timestamp 1662439860
transform -1 0 3496 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  x4_x81
timestamp 1662439860
transform 1 0 1564 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x82
timestamp 1662439860
transform -1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x4_x83_x1
timestamp 1662439860
transform 1 0 9752 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x83_x2
timestamp 1662439860
transform 1 0 9844 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x83_x3
timestamp 1662439860
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x4_x84_x1
timestamp 1662439860
transform 1 0 6164 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x84_x2
timestamp 1662439860
transform 1 0 5060 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x84_x3
timestamp 1662439860
transform 1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x4_x85_x1
timestamp 1662439860
transform -1 0 2944 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x4_x85_x2
timestamp 1662439860
transform 1 0 3036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x4_x85_x3
timestamp 1662439860
transform -1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x86
timestamp 1662439860
transform 1 0 9292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x87
timestamp 1662439860
transform 1 0 7636 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x88
timestamp 1662439860
transform -1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x89
timestamp 1662439860
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4_x90
timestamp 1662439860
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x91
timestamp 1662439860
transform 1 0 9108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x92
timestamp 1662439860
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x93
timestamp 1662439860
transform 1 0 3956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x94
timestamp 1662439860
transform 1 0 4508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x95
timestamp 1662439860
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x4_x96
timestamp 1662439860
transform 1 0 1564 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x4_x97
timestamp 1662439860
transform 1 0 2300 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x4_x98
timestamp 1662439860
transform 1 0 1748 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  x4_x99
timestamp 1662439860
transform -1 0 18584 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x100
timestamp 1662439860
transform 1 0 17112 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x4_x102
timestamp 1662439860
transform 1 0 18216 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x103
timestamp 1662439860
transform -1 0 18584 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x104
timestamp 1662439860
transform 1 0 17848 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x105
timestamp 1662439860
transform -1 0 17940 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x106
timestamp 1662439860
transform 1 0 15364 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x107
timestamp 1662439860
transform -1 0 16008 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x108
timestamp 1662439860
transform 1 0 12512 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x109
timestamp 1662439860
transform 1 0 13984 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x110
timestamp 1662439860
transform 1 0 11684 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x111
timestamp 1662439860
transform -1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x112
timestamp 1662439860
transform 1 0 11684 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x113
timestamp 1662439860
transform 1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x114
timestamp 1662439860
transform 1 0 10672 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x115
timestamp 1662439860
transform -1 0 12696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x116
timestamp 1662439860
transform 1 0 9292 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x117
timestamp 1662439860
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  x4_x118
timestamp 1662439860
transform 1 0 7912 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4_x119
timestamp 1662439860
transform 1 0 8096 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x4_x132
timestamp 1662439860
transform -1 0 3404 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x4_x133
timestamp 1662439860
transform -1 0 3312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x5_x1
timestamp 1662439860
transform -1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x5_x2
timestamp 1662439860
transform 1 0 2576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  x5_x3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 2576 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  x5_x4
timestamp 1662439860
transform -1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  x5_x5
timestamp 1662439860
transform -1 0 5060 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x5_x6
timestamp 1662439860
transform 1 0 1932 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  x5_x7
timestamp 1662439860
transform 1 0 2300 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x8
timestamp 1662439860
transform 1 0 3956 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x9
timestamp 1662439860
transform -1 0 5980 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x10
timestamp 1662439860
transform 1 0 5060 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x11
timestamp 1662439860
transform 1 0 6532 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x12
timestamp 1662439860
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x13
timestamp 1662439860
transform -1 0 8832 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x14
timestamp 1662439860
transform 1 0 9200 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x15
timestamp 1662439860
transform 1 0 10120 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x16
timestamp 1662439860
transform 1 0 11040 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x17
timestamp 1662439860
transform 1 0 11776 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x18
timestamp 1662439860
transform 1 0 13984 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x19
timestamp 1662439860
transform -1 0 16100 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x20
timestamp 1662439860
transform -1 0 6624 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  x5_x21
timestamp 1662439860
transform 1 0 5980 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_1  x5_x22
timestamp 1662439860
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x5_x23
timestamp 1662439860
transform -1 0 2576 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x5_x24
timestamp 1662439860
transform -1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x5_x25
timestamp 1662439860
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x5_x26
timestamp 1662439860
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x5_x27
timestamp 1662439860
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x5_x28
timestamp 1662439860
transform -1 0 2576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  x6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 17848 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x7_x1
timestamp 1662439860
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  x7_x2
timestamp 1662439860
transform -1 0 2300 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x7_x3
timestamp 1662439860
transform 1 0 1656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x7_x4
timestamp 1662439860
transform 1 0 3312 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x7_x5
timestamp 1662439860
transform 1 0 3956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x7_x6
timestamp 1662439860
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  x7_x9
timestamp 1662439860
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x7_x14
timestamp 1662439860
transform -1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  x7_x17
timestamp 1662439860
transform 1 0 2208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  x7_x19
timestamp 1662439860
transform -1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x7_x26
timestamp 1662439860
transform -1 0 5428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x7_x27
timestamp 1662439860
transform -1 0 5520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x25
timestamp 1662439860
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x26
timestamp 1662439860
transform -1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x27
timestamp 1662439860
transform -1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x28
timestamp 1662439860
transform 1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x29
timestamp 1662439860
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  x30
timestamp 1662439860
transform -1 0 18032 0 -1 10880
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 VDD
port 0 nsew signal bidirectional
flabel metal4 s 5842 2128 6162 21808 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 10741 2128 11061 21808 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 15640 2128 15960 21808 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 20539 2128 20859 21808 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 3393 2128 3713 21808 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 8292 2128 8612 21808 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 13191 2128 13511 21808 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 18090 2128 18410 21808 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 VSS
port 3 nsew signal bidirectional
flabel metal3 s 21061 17280 21861 17400 0 FreeSans 480 0 0 0 bit1
port 4 nsew signal tristate
flabel metal3 s 21061 1368 21861 1488 0 FreeSans 480 0 0 0 bit10
port 5 nsew signal tristate
flabel metal3 s 21061 15512 21861 15632 0 FreeSans 480 0 0 0 bit2
port 6 nsew signal tristate
flabel metal3 s 21061 13744 21861 13864 0 FreeSans 480 0 0 0 bit3
port 7 nsew signal tristate
flabel metal3 s 21061 11976 21861 12096 0 FreeSans 480 0 0 0 bit4
port 8 nsew signal tristate
flabel metal3 s 21061 10208 21861 10328 0 FreeSans 480 0 0 0 bit5
port 9 nsew signal tristate
flabel metal3 s 21061 8440 21861 8560 0 FreeSans 480 0 0 0 bit6
port 10 nsew signal tristate
flabel metal3 s 21061 6672 21861 6792 0 FreeSans 480 0 0 0 bit7
port 11 nsew signal tristate
flabel metal3 s 21061 4904 21861 5024 0 FreeSans 480 0 0 0 bit8
port 12 nsew signal tristate
flabel metal3 s 21061 3136 21861 3256 0 FreeSans 480 0 0 0 bit9
port 13 nsew signal tristate
flabel metal3 s 21061 20816 21861 20936 0 FreeSans 480 0 0 0 clk
port 14 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 comp_out_n
port 15 nsew signal input
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 comp_out_p
port 16 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 comparator_clk
port 17 nsew signal tristate
flabel metal3 s 21061 19048 21861 19168 0 FreeSans 480 0 0 0 done
port 18 nsew signal tristate
flabel metal3 s 21061 22584 21861 22704 0 FreeSans 480 0 0 0 reset
port 19 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 sw_n1
port 20 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 sw_n2
port 21 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 sw_n3
port 22 nsew signal tristate
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 sw_n4
port 23 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 sw_n5
port 24 nsew signal tristate
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 sw_n6
port 25 nsew signal tristate
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 sw_n7
port 26 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 sw_n8
port 27 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 sw_n_sp1
port 28 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 sw_n_sp2
port 29 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 sw_n_sp3
port 30 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 sw_n_sp4
port 31 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 sw_n_sp5
port 32 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 sw_n_sp6
port 33 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 sw_n_sp7
port 34 nsew signal tristate
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 sw_n_sp8
port 35 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 sw_n_sp9
port 36 nsew signal tristate
flabel metal2 s 18602 23205 18658 24005 0 FreeSans 224 90 0 0 sw_p1
port 37 nsew signal tristate
flabel metal2 s 17314 23205 17370 24005 0 FreeSans 224 90 0 0 sw_p2
port 38 nsew signal tristate
flabel metal2 s 12162 23205 12218 24005 0 FreeSans 224 90 0 0 sw_p3
port 39 nsew signal tristate
flabel metal2 s 10874 23205 10930 24005 0 FreeSans 224 90 0 0 sw_p4
port 40 nsew signal tristate
flabel metal2 s 9586 23205 9642 24005 0 FreeSans 224 90 0 0 sw_p5
port 41 nsew signal tristate
flabel metal2 s 4434 23205 4490 24005 0 FreeSans 224 90 0 0 sw_p6
port 42 nsew signal tristate
flabel metal2 s 3146 23205 3202 24005 0 FreeSans 224 90 0 0 sw_p7
port 43 nsew signal tristate
flabel metal2 s 1858 23205 1914 24005 0 FreeSans 224 90 0 0 sw_p8
port 44 nsew signal tristate
flabel metal2 s 21178 23205 21234 24005 0 FreeSans 224 90 0 0 sw_p_sp1
port 45 nsew signal tristate
flabel metal2 s 19890 23205 19946 24005 0 FreeSans 224 90 0 0 sw_p_sp2
port 46 nsew signal tristate
flabel metal2 s 16026 23205 16082 24005 0 FreeSans 224 90 0 0 sw_p_sp3
port 47 nsew signal tristate
flabel metal2 s 14738 23205 14794 24005 0 FreeSans 224 90 0 0 sw_p_sp4
port 48 nsew signal tristate
flabel metal2 s 13450 23205 13506 24005 0 FreeSans 224 90 0 0 sw_p_sp5
port 49 nsew signal tristate
flabel metal2 s 8298 23205 8354 24005 0 FreeSans 224 90 0 0 sw_p_sp6
port 50 nsew signal tristate
flabel metal2 s 7010 23205 7066 24005 0 FreeSans 224 90 0 0 sw_p_sp7
port 51 nsew signal tristate
flabel metal2 s 5722 23205 5778 24005 0 FreeSans 224 90 0 0 sw_p_sp8
port 52 nsew signal tristate
flabel metal2 s 570 23205 626 24005 0 FreeSans 224 90 0 0 sw_p_sp9
port 53 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 sw_sample
port 54 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 21861 24005
<< end >>
