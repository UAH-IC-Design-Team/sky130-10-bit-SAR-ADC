magic
tech sky130A
timestamp 1667663783
<< metal4 >>
rect 250 0 300 600
rect 600 0 650 600
rect 1050 0 1100 600
rect 1400 0 1450 600
rect 1850 0 1900 600
rect 2200 0 2250 600
rect 2650 0 2700 600
rect 3000 0 3050 600
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
array 0 3 800 0 0 800
timestamp 1667663783
transform 1 0 325 0 1 300
box -325 -300 325 300
<< end >>
