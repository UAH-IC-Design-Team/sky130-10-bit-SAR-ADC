magic
tech sky130A
magscale 1 2
timestamp 1667523134
<< nwell >>
rect 11420 8540 12410 8880
rect 10660 7540 13060 7880
rect 7730 6100 8510 6110
rect 7730 6080 8620 6100
rect 7731 5834 8620 6080
rect 8841 5900 9780 6110
rect 7730 5779 8620 5834
rect 8840 5779 9780 5900
rect 11060 5800 12680 7280
rect 14180 5780 16410 6110
rect 14190 5779 14442 5780
rect 14550 5779 14796 5780
rect 15190 5779 15432 5780
rect 7320 5080 10240 5410
rect 8110 5079 8356 5080
rect 8930 5079 9176 5080
rect 9750 5079 10398 5080
rect 7540 4370 10150 4710
<< nsubdiff >>
rect 11120 7070 11240 7100
rect 11120 6940 11240 6970
rect 12520 7070 12640 7100
rect 12520 6940 12640 6970
rect 11120 6830 11240 6860
rect 11120 6700 11240 6730
rect 12520 6830 12640 6860
rect 12520 6700 12640 6730
<< nsubdiffcont >>
rect 11120 6970 11240 7070
rect 12520 6970 12640 7070
rect 11120 6730 11240 6830
rect 12520 6730 12640 6830
<< locali >>
rect 11120 7070 11240 7090
rect 11120 6950 11240 6970
rect 12520 7070 12640 7090
rect 12520 6950 12640 6970
rect 11120 6830 11240 6850
rect 11120 6710 11240 6730
rect 12520 6830 12640 6850
rect 12520 6710 12640 6730
rect 8312 5733 8830 5773
rect 9106 5733 9340 5780
rect 14500 5733 14652 5781
rect 15000 5733 15490 5773
rect 8031 5029 8290 5083
rect 8851 5033 9105 5076
rect 9670 5013 9910 5090
rect 9670 5010 9679 5013
rect 7703 4315 7853 4389
rect 9760 4381 9807 4390
rect 8076 4337 8312 4381
rect 8670 4333 9148 4373
rect 9760 4329 9920 4381
rect 9760 4320 9807 4329
<< viali >>
rect 11120 6970 11240 7070
rect 12520 6970 12640 7070
rect 11120 6730 11240 6830
rect 12520 6730 12640 6830
rect 10037 5232 10071 5266
rect 10037 5158 10071 5192
rect 10038 4919 10072 4953
<< metal1 >>
rect 10700 7570 11150 7820
rect 10700 7130 11030 7570
rect 11550 7380 11670 7730
rect 11760 7620 11960 7780
rect 7458 6014 9740 6110
rect 9910 5870 10330 7020
rect 10470 6630 11030 7130
rect 11110 7270 11670 7380
rect 11110 7070 11250 7270
rect 11110 6970 11120 7070
rect 11240 6970 11250 7070
rect 11110 6830 11250 6970
rect 11110 6730 11120 6830
rect 11240 6730 11250 6830
rect 11110 6710 11250 6730
rect 10470 6520 11330 6630
rect 10470 6210 11030 6520
rect 10470 6110 11330 6210
rect 11380 5940 11510 7230
rect 11550 6890 11670 7270
rect 12080 7380 12200 7730
rect 12570 7570 12980 7820
rect 12080 7270 12650 7380
rect 11730 6770 11820 7190
rect 11930 7090 12020 7190
rect 11930 7020 11940 7090
rect 12010 7020 12020 7090
rect 11930 6910 12020 7020
rect 11930 6840 11940 6910
rect 12010 6840 12020 6910
rect 12080 6890 12200 7270
rect 11930 6810 12020 6840
rect 11730 6690 12200 6770
rect 11550 6670 11660 6680
rect 11550 6610 11590 6670
rect 11650 6610 11660 6670
rect 11550 6570 11660 6610
rect 11550 6510 11590 6570
rect 11650 6510 11660 6570
rect 11550 6470 11660 6510
rect 11550 6410 11590 6470
rect 11650 6410 11660 6470
rect 9910 5690 10740 5870
rect 11550 5810 11660 6410
rect 12090 5980 12200 6690
rect 12090 5900 12100 5980
rect 12190 5900 12200 5980
rect 12240 5940 12370 7230
rect 12510 7070 12650 7270
rect 12510 6970 12520 7070
rect 12640 6970 12650 7070
rect 12510 6830 12650 6970
rect 12510 6730 12520 6830
rect 12640 6730 12650 6830
rect 12510 6710 12650 6730
rect 12720 7120 12980 7570
rect 12720 6630 13260 7120
rect 12420 6530 13260 6630
rect 12720 6200 13260 6530
rect 12420 6100 13260 6200
rect 12090 5850 12200 5900
rect 13400 5870 13820 7020
rect 14088 6014 16370 6110
rect 11200 5800 12060 5810
rect 11200 5690 11210 5800
rect 11270 5690 11320 5800
rect 11380 5690 11430 5800
rect 11490 5740 12060 5800
rect 11490 5690 11660 5740
rect 7458 5470 9740 5570
rect 7350 5310 10360 5410
rect 10030 5266 10130 5280
rect 10030 5232 10037 5266
rect 10071 5232 10130 5266
rect 10030 5220 10130 5232
rect 10030 5192 10040 5220
rect 10030 5158 10037 5192
rect 10030 5140 10040 5158
rect 10120 5140 10130 5220
rect 10030 5100 10130 5140
rect 10030 5020 10040 5100
rect 10120 5020 10130 5100
rect 10030 4953 10130 5020
rect 10460 5180 10740 5690
rect 11050 5550 11160 5690
rect 11050 5470 11060 5550
rect 11150 5470 11160 5550
rect 11050 5450 11160 5470
rect 11050 5370 11060 5450
rect 11150 5370 11160 5450
rect 11050 5320 11160 5370
rect 11200 5680 11660 5690
rect 11200 5290 11260 5680
rect 11300 5390 11550 5630
rect 11590 5300 11660 5680
rect 11690 5660 11770 5700
rect 11690 5600 11700 5660
rect 11760 5600 11770 5660
rect 11690 5550 11770 5600
rect 11690 5490 11700 5550
rect 11760 5490 11770 5550
rect 11690 5330 11770 5490
rect 11980 5330 12060 5740
rect 12090 5770 12100 5850
rect 12190 5810 12200 5850
rect 12190 5770 12540 5810
rect 12090 5680 12540 5770
rect 12090 5290 12160 5680
rect 12200 5390 12450 5630
rect 12490 5290 12540 5680
rect 12590 5550 12700 5700
rect 12590 5470 12600 5550
rect 12690 5470 12700 5550
rect 12590 5450 12700 5470
rect 12590 5370 12600 5450
rect 12690 5370 12700 5450
rect 12590 5330 12700 5370
rect 12990 5690 13820 5870
rect 12990 5180 13270 5690
rect 14088 5470 16360 5570
rect 10460 5000 13270 5180
rect 10030 4919 10038 4953
rect 10072 4919 10130 4953
rect 10030 4900 10130 4919
rect 7350 4770 10360 4870
rect 7450 4610 10180 4710
rect 11540 4500 12280 5000
rect 12620 4360 13430 4840
rect 7450 4070 10180 4170
<< via1 >>
rect 11940 7020 12010 7090
rect 11940 6840 12010 6910
rect 11590 6610 11650 6670
rect 11590 6510 11650 6570
rect 11590 6410 11650 6470
rect 12100 5900 12190 5980
rect 11210 5690 11270 5800
rect 11320 5690 11380 5800
rect 11430 5690 11490 5800
rect 10040 5192 10120 5220
rect 10040 5158 10071 5192
rect 10071 5158 10120 5192
rect 10040 5140 10120 5158
rect 10040 5020 10120 5100
rect 11060 5470 11150 5550
rect 11060 5370 11150 5450
rect 11700 5600 11760 5660
rect 11700 5490 11760 5550
rect 12100 5770 12190 5850
rect 12600 5470 12690 5550
rect 12600 5370 12690 5450
<< metal2 >>
rect 11930 7090 12020 7120
rect 11930 7020 11940 7090
rect 12010 7020 12020 7090
rect 11930 6910 12020 7020
rect 11930 6840 11940 6910
rect 12010 6840 12020 6910
rect 11930 6770 12020 6840
rect 11580 6690 12020 6770
rect 11580 6670 11660 6690
rect 11580 6610 11590 6670
rect 11650 6610 11660 6670
rect 11580 6570 11660 6610
rect 11580 6510 11590 6570
rect 11650 6510 11660 6570
rect 11580 6470 11660 6510
rect 11580 6410 11590 6470
rect 11650 6410 11660 6470
rect 11580 6400 11660 6410
rect 12090 5980 12200 5990
rect 12090 5900 12100 5980
rect 12190 5900 12200 5980
rect 12090 5850 12200 5900
rect 12090 5810 12100 5850
rect 9470 5800 11550 5810
rect 9470 5690 11210 5800
rect 11270 5690 11320 5800
rect 11380 5690 11430 5800
rect 11490 5690 11550 5800
rect 9470 5680 11550 5690
rect 11690 5770 12100 5810
rect 12190 5810 12200 5850
rect 12190 5770 13850 5810
rect 11690 5740 13850 5770
rect 11690 5660 11770 5740
rect 12090 5680 13850 5740
rect 11690 5600 11700 5660
rect 11760 5600 11770 5660
rect 11050 5550 11160 5560
rect 11050 5470 11060 5550
rect 11150 5470 11160 5550
rect 11690 5550 11770 5600
rect 11690 5490 11700 5550
rect 11760 5490 11770 5550
rect 11690 5480 11770 5490
rect 12590 5550 12700 5560
rect 11050 5460 11160 5470
rect 10030 5450 11160 5460
rect 12590 5470 12600 5550
rect 12690 5470 12700 5550
rect 12590 5450 12700 5470
rect 10030 5370 11060 5450
rect 11150 5370 12600 5450
rect 12690 5370 12700 5450
rect 10030 5360 12700 5370
rect 10030 5220 10130 5360
rect 10030 5140 10040 5220
rect 10120 5140 10130 5220
rect 10030 5100 10130 5140
rect 10030 5020 10040 5100
rect 10120 5020 10130 5100
rect 10030 5010 10130 5020
use sky130_fd_pr__pfet_01v8_FBQ47L  XM1
timestamp 1666924120
transform 0 1 12500 1 0 7701
box -161 -600 169 560
use sky130_fd_pr__pfet_01v8_5AQ4BN  XM2
timestamp 1666923623
transform 0 -1 11220 1 0 7701
box -161 -620 179 560
use sky130_fd_pr__nfet_01v8_ZRN2GS  XM4
timestamp 1667435063
transform 0 -1 10398 -1 0 6609
box -509 -532 509 598
use sky130_fd_pr__nfet_01v8_ZCCU26  XM9
timestamp 1667500205
transform 0 1 12448 -1 0 4669
box -269 -1088 269 1028
use sky130_fd_pr__nfet_01v8_ZZU2YL  XM13
timestamp 1667436771
transform 0 1 11279 -1 0 5511
box -221 -179 221 119
use sky130_fd_pr__nfet_01v8_ZRN2GS  sky130_fd_pr__nfet_01v8_ZRN2GS_0
timestamp 1667435063
transform 0 1 13332 1 0 6609
box -509 -532 509 598
use sky130_fd_pr__nfet_01v8_ZZU2YL  sky130_fd_pr__nfet_01v8_ZZU2YL_0
timestamp 1667436771
transform 0 1 12179 1 0 5511
box -221 -179 221 119
use sky130_fd_pr__nfet_01v8_ZZU2YL  sky130_fd_pr__nfet_01v8_ZZU2YL_1
timestamp 1667436771
transform 0 -1 11569 1 0 5511
box -221 -179 221 119
use sky130_fd_pr__nfet_01v8_ZZU2YL  sky130_fd_pr__nfet_01v8_ZZU2YL_2
timestamp 1667436771
transform 0 -1 12469 1 0 5511
box -221 -179 221 119
use sky130_fd_pr__pfet_01v8_QPTUVJ  sky130_fd_pr__pfet_01v8_QPTUVJ_0
timestamp 1667435677
transform 0 -1 11529 1 0 7007
box -257 -271 263 219
use sky130_fd_pr__pfet_01v8_QPTUVJ  sky130_fd_pr__pfet_01v8_QPTUVJ_1
timestamp 1667435677
transform 0 1 12221 1 0 7007
box -257 -271 263 219
use sky130_fd_pr__pfet_01v8_RPBXXN  sky130_fd_pr__pfet_01v8_RPBXXN_0
timestamp 1666924247
transform 0 -1 12221 -1 0 6249
box -451 -269 449 221
use sky130_fd_pr__pfet_01v8_RPBXXN  sky130_fd_pr__pfet_01v8_RPBXXN_1
timestamp 1666924247
transform 0 1 11529 -1 0 6249
box -451 -269 449 221
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 10268 0 1 4818
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1662439860
transform 1 0 14088 0 1 5518
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1662439860
transform 1 0 9648 0 1 5518
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1662439860
transform 1 0 10088 0 1 4118
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  x1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14258 0 1 5518
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14618 0 1 5518
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 15258 0 1 5518
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x4
timestamp 1662439860
transform -1 0 9564 0 1 5518
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x5
timestamp 1662439860
transform -1 0 9200 0 1 5518
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x6
timestamp 1662439860
transform -1 0 8562 0 1 5518
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x7
timestamp 1662439860
transform 1 0 7458 0 1 4118
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 7358 0 1 4818
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9818 0 1 4818
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x10
timestamp 1662439860
transform 1 0 8178 0 1 4818
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8998 0 1 4818
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x12
timestamp 1662439860
transform 1 0 7818 0 1 4118
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  x13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 11458 0 1 8288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x14
timestamp 1662439860
transform 1 0 8268 0 1 4118
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x15
timestamp 1662439860
transform 1 0 8898 0 1 4118
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  x16
timestamp 1662439860
transform 1 0 11818 0 1 8288
box -38 -48 590 592
<< labels >>
flabel nwell s 8518 6045 8552 6079 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
<< end >>
