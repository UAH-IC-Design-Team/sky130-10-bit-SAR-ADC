magic
tech sky130A
magscale 1 2
timestamp 1665684523
<< metal1 >>
rect -74500 56680 -74300 56880
rect -82840 56180 -82640 56380
rect -96720 55840 -96520 56040
rect -64300 55980 -64100 56180
rect -59520 56020 -59320 56220
rect -57440 55760 -57240 55960
rect -55920 55900 -55720 56100
rect -54080 56000 -53880 56200
rect -49940 56000 -49740 56200
rect -51560 55680 -51360 55880
rect -47860 24000 -47660 24200
rect -45360 23880 -45160 24080
rect -44040 23900 -43840 24100
rect -42180 23820 -41980 24020
rect -39540 23820 -39340 24020
rect -38100 23700 -37900 23900
rect -37160 23660 -36960 23860
rect -36640 18660 -36440 18860
rect -36640 18220 -36440 18420
rect -47940 13040 -47740 13240
rect -45440 13020 -45240 13220
rect -44020 12980 -43820 13180
rect -41540 13120 -41340 13320
rect -39260 13160 -39060 13360
rect -38160 13200 -37960 13400
rect -37140 13120 -36940 13320
rect -92280 -18800 -92080 -18600
rect -73400 -19040 -73200 -18840
rect -57440 -18900 -57240 -18700
rect -56000 -18800 -55800 -18600
rect -51340 -18920 -51140 -18720
rect -49900 -18920 -49700 -18720
rect -82880 -19300 -82680 -19100
rect -64640 -19320 -64440 -19120
rect -59920 -19220 -59720 -19020
rect -53880 -19180 -53680 -18980
<< metal3 >>
rect -97300 19000 -85816 55080
rect -85400 19000 -79668 55080
rect -79300 19000 -67816 55080
rect -67400 19000 -61668 55080
rect -61200 19000 -58344 55080
rect -58000 19000 -56582 55080
rect -56200 19000 -55501 55080
rect -55200 19000 -52344 55080
rect -52000 19000 -50582 55080
rect -50200 19000 -49501 55080
rect -49200 19000 -46344 23410
rect -46000 19000 -44582 23410
rect -44300 19000 -43601 23410
rect -43300 19000 -40444 23410
rect -40100 19000 -38682 23410
rect -38400 19000 -37701 23410
rect -37400 19000 -36701 23410
rect -97300 -18000 -85816 18080
rect -85400 -18000 -79668 18080
rect -79300 -18000 -67816 18080
rect -67400 -18000 -61668 18080
rect -61200 -18000 -58344 18080
rect -58000 -18000 -56582 18080
rect -56200 -18000 -55501 18080
rect -55200 -18000 -52344 18080
rect -52000 -18000 -50582 18080
rect -50200 -18000 -49501 18080
rect -49200 13700 -46344 18110
rect -46000 13700 -44582 18110
rect -44300 13700 -43601 18110
rect -43300 13700 -40444 18110
rect -40100 13700 -38682 18110
rect -38400 13700 -37701 18110
rect -37400 13700 -36701 18110
<< metal4 >>
rect -97060 55200 -86160 55300
rect -97060 55080 -96940 55200
rect -96340 55080 -96220 55200
rect -95620 55080 -95500 55200
rect -94900 55080 -94780 55200
rect -94180 55080 -94060 55200
rect -93460 55080 -93340 55200
rect -92740 55080 -92620 55200
rect -92020 55080 -91900 55200
rect -91300 55080 -91180 55200
rect -90580 55080 -90460 55200
rect -89860 55080 -89740 55200
rect -89160 55080 -89040 55200
rect -88440 55080 -88320 55200
rect -87720 55080 -87600 55200
rect -87000 55080 -86880 55200
rect -86280 55080 -86160 55200
rect -85160 55200 -80000 55300
rect -85160 55080 -85040 55200
rect -84440 55080 -84320 55200
rect -83720 55080 -83600 55200
rect -83000 55080 -82880 55200
rect -82280 55080 -82160 55200
rect -81560 55080 -81440 55200
rect -80840 55080 -80720 55200
rect -80120 55080 -80000 55200
rect -79060 55180 -68160 55280
rect -79060 55080 -78940 55180
rect -78340 55080 -78220 55180
rect -77620 55080 -77500 55180
rect -76900 55080 -76780 55180
rect -76180 55080 -76060 55180
rect -75460 55080 -75340 55180
rect -74740 55080 -74620 55180
rect -74020 55080 -73900 55180
rect -73300 55080 -73180 55180
rect -72580 55080 -72460 55180
rect -71860 55080 -71740 55180
rect -71160 55080 -71040 55180
rect -70440 55080 -70320 55180
rect -69720 55080 -69600 55180
rect -69000 55080 -68880 55180
rect -68280 55080 -68160 55180
rect -67060 55200 -61900 55300
rect -67060 55080 -66940 55200
rect -66340 55080 -66220 55200
rect -65620 55080 -65500 55200
rect -64900 55080 -64780 55200
rect -64180 55080 -64060 55200
rect -63460 55080 -63340 55200
rect -62740 55080 -62620 55200
rect -62020 55080 -61900 55200
rect -60960 55200 -58680 55300
rect -60960 55080 -60840 55200
rect -60240 55080 -60120 55200
rect -59520 55080 -59400 55200
rect -58800 55080 -58680 55200
rect -57760 55200 -56920 55300
rect -57760 55080 -57640 55200
rect -57040 55080 -56920 55200
rect -55960 55080 -55840 55300
rect -54960 55200 -52680 55300
rect -54960 55080 -54840 55200
rect -54240 55080 -54120 55200
rect -53520 55080 -53400 55200
rect -52800 55080 -52680 55200
rect -51760 55200 -50920 55300
rect -51760 55080 -51640 55200
rect -51040 55080 -50920 55200
rect -49960 55080 -49840 55300
rect -48980 23560 -46660 23700
rect -48980 23260 -48820 23560
rect -48260 23260 -48100 23560
rect -47540 23260 -47380 23560
rect -46820 23260 -46660 23560
rect -45780 23560 -44880 23680
rect -43080 23560 -40760 23680
rect -39880 23560 -39000 23680
rect -45780 23260 -45620 23560
rect -45040 23260 -44880 23560
rect -44080 23260 -43920 23560
rect -43080 23260 -42920 23560
rect -42360 23260 -42200 23560
rect -41640 23260 -41480 23560
rect -40920 23260 -40760 23560
rect -39860 23260 -39700 23560
rect -39160 23260 -39000 23560
rect -38180 23260 -38020 23560
rect -37180 23260 -37020 23560
rect -96740 18880 -96620 19000
rect -96020 18880 -95900 19000
rect -95300 18880 -95180 19000
rect -94580 18880 -94460 19000
rect -93860 18880 -93740 19000
rect -93140 18880 -93020 19000
rect -92420 18880 -92300 19000
rect -91700 18880 -91580 19000
rect -90980 18880 -90860 19000
rect -90260 18880 -90140 19000
rect -89540 18880 -89420 19000
rect -88840 18880 -88720 19000
rect -88120 18880 -88000 19000
rect -87400 18880 -87280 19000
rect -86680 18880 -86560 19000
rect -85960 18880 -85840 19000
rect -84840 18880 -84720 19000
rect -84120 18880 -84000 19000
rect -83400 18880 -83280 19000
rect -82680 18880 -82560 19000
rect -81960 18880 -81840 19000
rect -81240 18880 -81120 19000
rect -80520 18880 -80400 19000
rect -79800 18880 -79680 19000
rect -78740 18900 -78620 19000
rect -78020 18900 -77900 19000
rect -77300 18900 -77180 19000
rect -76580 18900 -76460 19000
rect -75860 18900 -75740 19000
rect -75140 18900 -75020 19000
rect -74420 18900 -74300 19000
rect -73700 18900 -73580 19000
rect -72980 18900 -72860 19000
rect -72260 18900 -72140 19000
rect -71540 18900 -71420 19000
rect -70840 18900 -70720 19000
rect -70120 18900 -70000 19000
rect -69400 18900 -69280 19000
rect -68680 18900 -68560 19000
rect -67960 18900 -67840 19000
rect -66740 18900 -66620 19000
rect -78740 18880 -66620 18900
rect -66020 18880 -65900 19000
rect -65300 18880 -65180 19000
rect -64580 18880 -64460 19000
rect -63860 18880 -63740 19000
rect -63140 18880 -63020 19000
rect -62420 18880 -62300 19000
rect -61700 18880 -61580 19000
rect -60640 18880 -60520 19000
rect -59920 18880 -59800 19000
rect -59200 18880 -59080 19000
rect -58480 18880 -58360 19000
rect -57440 18880 -57320 19000
rect -56720 18880 -56600 19000
rect -55640 18880 -55520 19000
rect -54640 18880 -54520 19000
rect -53920 18880 -53800 19000
rect -53200 18880 -53080 19000
rect -52480 18880 -52360 19000
rect -51440 18880 -51320 19000
rect -50720 18880 -50600 19000
rect -49640 18880 -49520 19000
rect -48600 18880 -48500 19020
rect -47880 18880 -47780 19020
rect -47160 18880 -47040 19020
rect -46460 18880 -46340 19020
rect -45420 18880 -45300 19020
rect -44700 18880 -44580 19020
rect -43720 18880 -43600 19020
rect -42720 18880 -42600 19020
rect -42000 18880 -41880 19020
rect -41280 18880 -41160 19020
rect -40560 18880 -40440 19020
rect -39520 18880 -39400 19020
rect -38800 18880 -38680 19020
rect -37800 18880 -37680 19020
rect -36800 18880 -36680 19020
rect -96740 18660 -36680 18880
rect -96740 18200 -36680 18420
rect -96740 18080 -96620 18200
rect -96020 18080 -95900 18200
rect -95300 18080 -95180 18200
rect -94580 18080 -94460 18200
rect -93860 18080 -93740 18200
rect -93140 18080 -93020 18200
rect -92420 18080 -92300 18200
rect -91700 18080 -91580 18200
rect -90980 18080 -90860 18200
rect -90260 18080 -90140 18200
rect -89540 18080 -89420 18200
rect -88840 18080 -88720 18200
rect -88120 18080 -88000 18200
rect -87400 18080 -87280 18200
rect -86680 18080 -86560 18200
rect -85960 18080 -85840 18200
rect -84840 18080 -84720 18200
rect -84120 18080 -84000 18200
rect -83400 18080 -83280 18200
rect -82680 18080 -82560 18200
rect -81960 18080 -81840 18200
rect -81240 18080 -81120 18200
rect -80520 18080 -80400 18200
rect -79800 18080 -79680 18200
rect -78740 18180 -66620 18200
rect -78740 18080 -78620 18180
rect -78020 18080 -77900 18180
rect -77300 18080 -77180 18180
rect -76580 18080 -76460 18180
rect -75860 18080 -75740 18180
rect -75140 18080 -75020 18180
rect -74420 18080 -74300 18180
rect -73700 18080 -73580 18180
rect -72980 18080 -72860 18180
rect -72260 18080 -72140 18180
rect -71540 18080 -71420 18180
rect -70840 18080 -70720 18180
rect -70120 18080 -70000 18180
rect -69400 18080 -69280 18180
rect -68680 18080 -68560 18180
rect -67960 18080 -67840 18180
rect -66740 18080 -66620 18180
rect -66020 18080 -65900 18200
rect -65300 18080 -65180 18200
rect -64580 18080 -64460 18200
rect -63860 18080 -63740 18200
rect -63140 18080 -63020 18200
rect -62420 18080 -62300 18200
rect -61700 18080 -61580 18200
rect -60640 18080 -60520 18200
rect -59920 18080 -59800 18200
rect -59200 18080 -59080 18200
rect -58480 18080 -58360 18200
rect -57440 18080 -57320 18200
rect -56720 18080 -56600 18200
rect -55640 18080 -55520 18200
rect -54640 18080 -54520 18200
rect -53920 18080 -53800 18200
rect -53200 18080 -53080 18200
rect -52480 18080 -52360 18200
rect -51440 18080 -51320 18200
rect -50720 18080 -50600 18200
rect -49640 18080 -49520 18200
rect -48600 18080 -48480 18200
rect -47880 18080 -47760 18200
rect -47160 18080 -47040 18200
rect -46440 18080 -46340 18200
rect -45400 18080 -45280 18200
rect -44680 18080 -44560 18200
rect -43700 18080 -43600 18200
rect -42700 18080 -42600 18200
rect -42000 18080 -41880 18200
rect -41280 18080 -41160 18200
rect -40560 18080 -40440 18200
rect -39520 18080 -39400 18200
rect -38800 18080 -38680 18200
rect -37820 18080 -37700 18200
rect -36820 18080 -36680 18200
rect -48980 13580 -48820 13840
rect -48260 13580 -48100 13840
rect -47540 13580 -47380 13840
rect -46820 13580 -46660 13840
rect -48980 13420 -46660 13580
rect -45780 13580 -45620 13840
rect -45060 13580 -44900 13840
rect -44080 13580 -43920 13840
rect -43080 13580 -42920 13840
rect -42360 13580 -42200 13840
rect -41660 13580 -41500 13840
rect -40920 13580 -40760 13840
rect -45780 13420 -44900 13580
rect -43080 13420 -40760 13580
rect -39880 13580 -39720 13840
rect -39160 13580 -39000 13840
rect -38180 13580 -38020 13840
rect -37180 13580 -37020 13840
rect -39880 13420 -39000 13580
rect -97060 -18120 -96940 -18000
rect -96340 -18120 -96220 -18000
rect -95620 -18120 -95500 -18000
rect -94900 -18120 -94780 -18000
rect -94180 -18120 -94060 -18000
rect -93460 -18120 -93340 -18000
rect -92740 -18120 -92620 -18000
rect -92020 -18120 -91900 -18000
rect -91300 -18120 -91180 -18000
rect -90580 -18120 -90460 -18000
rect -89860 -18120 -89740 -18000
rect -89160 -18120 -89040 -18000
rect -88440 -18120 -88320 -18000
rect -87720 -18120 -87600 -18000
rect -87000 -18120 -86880 -18000
rect -86280 -18120 -86160 -18000
rect -97060 -18220 -86160 -18120
rect -85160 -18120 -85040 -18000
rect -84440 -18120 -84320 -18000
rect -83720 -18120 -83600 -18000
rect -83000 -18120 -82880 -18000
rect -82280 -18120 -82160 -18000
rect -81560 -18120 -81440 -18000
rect -80840 -18120 -80720 -18000
rect -80120 -18120 -80000 -18000
rect -85160 -18220 -80000 -18120
rect -79060 -18100 -78940 -18000
rect -78340 -18100 -78220 -18000
rect -77620 -18100 -77500 -18000
rect -76900 -18100 -76780 -18000
rect -76180 -18100 -76060 -18000
rect -75460 -18100 -75340 -18000
rect -74740 -18100 -74620 -18000
rect -74020 -18100 -73900 -18000
rect -73300 -18100 -73180 -18000
rect -72580 -18100 -72460 -18000
rect -71860 -18100 -71740 -18000
rect -71160 -18100 -71040 -18000
rect -70440 -18100 -70320 -18000
rect -69720 -18100 -69600 -18000
rect -69000 -18100 -68880 -18000
rect -68280 -18100 -68160 -18000
rect -79060 -18200 -68160 -18100
rect -67060 -18120 -66940 -18000
rect -66340 -18120 -66220 -18000
rect -65620 -18120 -65500 -18000
rect -64900 -18120 -64780 -18000
rect -64180 -18120 -64060 -18000
rect -63460 -18120 -63340 -18000
rect -62740 -18120 -62620 -18000
rect -62020 -18120 -61900 -18000
rect -67060 -18220 -61900 -18120
rect -60960 -18120 -60840 -18000
rect -60240 -18120 -60120 -18000
rect -59520 -18120 -59400 -18000
rect -58800 -18120 -58680 -18000
rect -60960 -18220 -58680 -18120
rect -57760 -18120 -57640 -18000
rect -57040 -18120 -56920 -18000
rect -57760 -18220 -56920 -18120
rect -55960 -18220 -55840 -18000
rect -54960 -18120 -54840 -18000
rect -54240 -18120 -54120 -18000
rect -53520 -18120 -53400 -18000
rect -52800 -18120 -52680 -18000
rect -54960 -18220 -52680 -18120
rect -51760 -18120 -51640 -18000
rect -51040 -18120 -50920 -18000
rect -51760 -18220 -50920 -18120
rect -49960 -18220 -49840 -18000
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  XC1
timestamp 1665161463
transform 1 0 -73558 0 1 37040
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  XC2
timestamp 1665159686
transform 1 0 -64434 0 1 40
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  XC4
timestamp 1665159686
transform 1 0 -82534 0 1 40
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  XC5
timestamp 1665159686
transform 1 0 -53772 0 1 40
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  XC6
timestamp 1665159686
transform 1 0 -57291 0 1 37040
box -709 -18040 709 18040
use sky130_fd_pr__cap_mim_m3_1_LSQHR5  XC7
timestamp 1665159686
transform 1 0 -55850 0 1 37040
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  XC8
timestamp 1665159686
transform 1 0 -53772 0 1 37040
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  XC9
timestamp 1665159686
transform 1 0 -51291 0 1 37040
box -709 -18040 709 18040
use sky130_fd_pr__cap_mim_m3_1_EDBB5V  XC10
timestamp 1665159686
transform 1 0 -49850 0 1 37040
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_LQ5JR5  XC11
timestamp 1665675118
transform 1 0 -47772 0 1 15905
box -1428 -2205 1428 2205
use sky130_fd_pr__cap_mim_m3_1_LQPHR5  XC12
timestamp 1665675118
transform 1 0 -39391 0 1 21205
box -709 -2205 709 2205
use sky130_fd_pr__cap_mim_m3_1_EXCB5V  XC13
timestamp 1665159686
transform 1 0 -37050 0 1 15905
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_EXCB5V  XC16
timestamp 1665159686
transform 1 0 -37050 0 1 21205
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_EXCB5V  XC17
timestamp 1665159686
transform 1 0 -38050 0 1 15905
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  XC18
timestamp 1665161463
transform 1 0 -91558 0 1 37040
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  XC19
timestamp 1665159686
transform 1 0 -64434 0 1 37040
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  XC23
timestamp 1665159686
transform 1 0 -51291 0 1 40
box -709 -18040 709 18040
use sky130_fd_pr__cap_mim_m3_1_EDBB5V  XC24
timestamp 1665159686
transform 1 0 -55850 0 1 40
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_LSQHR5  XC27
timestamp 1665159686
transform 1 0 -49850 0 1 40
box -350 -18040 349 18040
use sky130_fd_pr__cap_mim_m3_1_LQ5JR5  XC28
timestamp 1665675118
transform 1 0 -41872 0 1 21205
box -1428 -2205 1428 2205
use sky130_fd_pr__cap_mim_m3_1_LQPHR5  XC29
timestamp 1665675118
transform 1 0 -45291 0 1 15905
box -709 -2205 709 2205
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  XC30
timestamp 1665161463
transform 1 0 -38050 0 1 21205
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_LQ5JR5  XC31
timestamp 1665675118
transform 1 0 -47772 0 1 21205
box -1428 -2205 1428 2205
use sky130_fd_pr__cap_mim_m3_1_LQPHR5  XC32
timestamp 1665675118
transform 1 0 -45291 0 1 21205
box -709 -2205 709 2205
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  XC33
timestamp 1665161463
transform 1 0 -43950 0 1 15905
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_LQSHR5  XC34
timestamp 1665161463
transform 1 0 -43950 0 1 21205
box -350 -2205 349 2205
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  sky130_fd_pr__cap_mim_m3_1_9SQ6B5_0
timestamp 1665161463
transform 1 0 -91558 0 1 40
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_9SQ6B5  sky130_fd_pr__cap_mim_m3_1_9SQ6B5_1
timestamp 1665161463
transform 1 0 -73558 0 1 40
box -5742 -18040 5742 18040
use sky130_fd_pr__cap_mim_m3_1_LQ5JR5  sky130_fd_pr__cap_mim_m3_1_LQ5JR5_0
timestamp 1665675118
transform 1 0 -41872 0 1 15905
box -1428 -2205 1428 2205
use sky130_fd_pr__cap_mim_m3_1_LQPHR5  sky130_fd_pr__cap_mim_m3_1_LQPHR5_0
timestamp 1665675118
transform 1 0 -39391 0 1 15905
box -709 -2205 709 2205
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  sky130_fd_pr__cap_mim_m3_1_LS3JR5_0
timestamp 1665159686
transform 1 0 -59772 0 1 40
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LS3JR5  sky130_fd_pr__cap_mim_m3_1_LS3JR5_1
timestamp 1665159686
transform 1 0 -59772 0 1 37040
box -1428 -18040 1428 18040
use sky130_fd_pr__cap_mim_m3_1_LSFHR5  sky130_fd_pr__cap_mim_m3_1_LSFHR5_0
timestamp 1665159686
transform 1 0 -82534 0 1 37040
box -2866 -18040 2866 18040
use sky130_fd_pr__cap_mim_m3_1_LSVHR5  sky130_fd_pr__cap_mim_m3_1_LSVHR5_0
timestamp 1665159686
transform 1 0 -57291 0 1 40
box -709 -18040 709 18040
<< labels >>
flabel metal1 -36640 18220 -36440 18420 0 FreeSans 256 0 0 0 Vin_n
port 11 nsew
flabel metal1 -37140 13120 -36940 13320 0 FreeSans 256 0 0 0 sw_sp_n9
port 0 nsew
flabel metal1 -44020 12980 -43820 13180 0 FreeSans 256 0 0 0 sw_sp_n8
port 1 nsew
flabel metal1 -45440 13020 -45240 13220 0 FreeSans 256 0 0 0 sw_sp_n7
port 2 nsew
flabel metal1 -47940 13040 -47740 13240 0 FreeSans 256 0 0 0 sw_sp_n6
port 3 nsew
flabel metal1 -56000 -18800 -55800 -18600 0 FreeSans 256 0 0 0 sw_sp_n5
port 4 nsew
flabel metal1 -57440 -18900 -57240 -18700 0 FreeSans 256 0 0 0 sw_sp_n4
port 5 nsew
flabel metal1 -59920 -19220 -59720 -19020 0 FreeSans 256 0 0 0 sw_sp_n3
port 6 nsew
flabel metal1 -82880 -19300 -82680 -19100 0 FreeSans 256 0 0 0 sw_sp_n2
port 7 nsew
flabel metal1 -92280 -18800 -92080 -18600 0 FreeSans 256 0 0 0 sw_sp_n1
port 9 nsew
flabel metal1 -37160 23660 -36960 23860 0 FreeSans 256 0 0 0 sw_sp_p9
port 12 nsew
flabel metal1 -44040 23900 -43840 24100 0 FreeSans 256 0 0 0 sw_sp_p8
port 13 nsew
flabel metal1 -45360 23880 -45160 24080 0 FreeSans 256 0 0 0 sw_sp_p7
port 14 nsew
flabel metal1 -47860 24000 -47660 24200 0 FreeSans 256 0 0 0 sw_sp_p6
port 15 nsew
flabel metal1 -55920 55900 -55720 56100 0 FreeSans 256 0 0 0 sw_sp_p5
port 16 nsew
flabel metal1 -57440 55760 -57240 55960 0 FreeSans 256 0 0 0 sw_sp_p4
port 17 nsew
flabel metal1 -59520 56020 -59320 56220 0 FreeSans 256 0 0 0 sw_sp_p3
port 18 nsew
flabel metal1 -82840 56180 -82640 56380 0 FreeSans 256 0 0 0 sw_sp_p2
port 19 nsew
flabel metal1 -38100 23700 -37900 23900 0 FreeSans 256 0 0 0 sw_p8
port 21 nsew
flabel metal1 -39540 23820 -39340 24020 0 FreeSans 256 0 0 0 sw_p7
port 23 nsew
flabel metal1 -42180 23820 -41980 24020 0 FreeSans 256 0 0 0 sw_p6
port 24 nsew
flabel metal1 -49940 56000 -49740 56200 0 FreeSans 256 0 0 0 sw_p5
port 25 nsew
flabel metal1 -51560 55680 -51360 55880 0 FreeSans 256 0 0 0 sw_p4
port 26 nsew
flabel metal1 -54080 56000 -53880 56200 0 FreeSans 256 0 0 0 sw_p3
port 27 nsew
flabel metal1 -64300 55980 -64100 56180 0 FreeSans 256 0 0 0 sw_p2
port 28 nsew
flabel metal1 -74500 56680 -74300 56880 0 FreeSans 256 0 0 0 sw_p1
port 29 nsew
flabel metal1 -38160 13200 -37960 13400 0 FreeSans 256 0 0 0 sw_n8
port 30 nsew
flabel metal1 -39260 13160 -39060 13360 0 FreeSans 256 0 0 0 sw_n7
port 31 nsew
flabel metal1 -41540 13120 -41340 13320 0 FreeSans 256 0 0 0 sw_n6
port 32 nsew
flabel metal1 -49900 -18920 -49700 -18720 0 FreeSans 256 0 0 0 sw_n5
port 33 nsew
flabel metal1 -51340 -18920 -51140 -18720 0 FreeSans 256 0 0 0 sw_n4
port 34 nsew
flabel metal1 -53880 -19180 -53680 -18980 0 FreeSans 256 0 0 0 sw_n3
port 35 nsew
flabel metal1 -64640 -19320 -64440 -19120 0 FreeSans 256 0 0 0 sw_n2
port 36 nsew
flabel metal1 -73400 -19040 -73200 -18840 0 FreeSans 256 0 0 0 sw_n1
port 37 nsew
flabel metal1 -96720 55840 -96520 56040 0 FreeSans 256 0 0 0 sw_sp_p1
port 20 nsew
flabel metal1 -36640 18660 -36440 18860 0 FreeSans 256 0 0 0 Vin_p
port 10 nsew
<< end >>
