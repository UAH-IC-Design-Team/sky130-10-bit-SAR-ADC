** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/tests/demux2/demux2_test.sch
**.subckt demux2_test
V3 VDD GND 1.8V
V4 VSS GND 0
x1 select VDD VSS out_0 v_in out_1 demux2
V1 select GND PULSE 0 1.8V 0 1ns 1ns 10us 20us
V2 v_in GND PULSE 0 1.8V 0 1ns 1ns 7us 15us
**** begin user architecture code
 .lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


.options acct list
.temp 25
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
.control
tran 0.1u 100u
plot select v_in+2 out_0+4 out_1+6
write pulse_generator_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  src/demux2/demux2.sym # of pins=6
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sch
.subckt demux2  S VDD VSS OUT_0 IN OUT_1
*.ipin S
*.opin OUT_0
*.ipin IN
*.opin OUT_1
*.iopin VDD
*.iopin VSS
x1 net1 IN VSS VSS VDD VDD OUT_0 sky130_fd_sc_hd__and2_0
x2 S IN VSS VSS VDD VDD OUT_1 sky130_fd_sc_hd__and2_0
x3 S VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_1
.ends

.GLOBAL GND
.end
