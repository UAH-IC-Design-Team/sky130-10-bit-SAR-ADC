magic
tech sky130A
timestamp 1666638196
<< metal1 >>
rect 0 0 70000 70000
rect 70411 -93 140411 69907
<< end >>
