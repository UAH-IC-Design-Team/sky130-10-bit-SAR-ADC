* Simulating the demuxer.
* Include the Sky130 libraries
.lib "/foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.include "/foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice"

* Include the magic export
.include "./demux2.spice"

* instantiate the demux
Xdemux VPWR VGND S IN OUT_0 OUT_1 demux2

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin IN VGND pulse(0 1.8 1p 10p 10p 1n 2n)
Vsel S VGND pulse(0 1.8 1p 10p 10p 2n 5n)
.tran 10e-12 7e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot IN S+2 OUT_0+4 OUT_1+6
.endc

.end
