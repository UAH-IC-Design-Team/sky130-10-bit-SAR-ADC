magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -386 36092 386 36120
rect -386 31858 302 36092
rect 366 31858 386 36092
rect -386 31830 386 31858
rect -386 31562 386 31590
rect -386 27328 302 31562
rect 366 27328 386 31562
rect -386 27300 386 27328
rect -386 27032 386 27060
rect -386 22798 302 27032
rect 366 22798 386 27032
rect -386 22770 386 22798
rect -386 22502 386 22530
rect -386 18268 302 22502
rect 366 18268 386 22502
rect -386 18240 386 18268
rect -386 17972 386 18000
rect -386 13738 302 17972
rect 366 13738 386 17972
rect -386 13710 386 13738
rect -386 13442 386 13470
rect -386 9208 302 13442
rect 366 9208 386 13442
rect -386 9180 386 9208
rect -386 8912 386 8940
rect -386 4678 302 8912
rect 366 4678 386 8912
rect -386 4650 386 4678
rect -386 4382 386 4410
rect -386 148 302 4382
rect 366 148 386 4382
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -4382 302 -148
rect 366 -4382 386 -148
rect -386 -4410 386 -4382
rect -386 -4678 386 -4650
rect -386 -8912 302 -4678
rect 366 -8912 386 -4678
rect -386 -8940 386 -8912
rect -386 -9208 386 -9180
rect -386 -13442 302 -9208
rect 366 -13442 386 -9208
rect -386 -13470 386 -13442
rect -386 -13738 386 -13710
rect -386 -17972 302 -13738
rect 366 -17972 386 -13738
rect -386 -18000 386 -17972
rect -386 -18268 386 -18240
rect -386 -22502 302 -18268
rect 366 -22502 386 -18268
rect -386 -22530 386 -22502
rect -386 -22798 386 -22770
rect -386 -27032 302 -22798
rect 366 -27032 386 -22798
rect -386 -27060 386 -27032
rect -386 -27328 386 -27300
rect -386 -31562 302 -27328
rect 366 -31562 386 -27328
rect -386 -31590 386 -31562
rect -386 -31858 386 -31830
rect -386 -36092 302 -31858
rect 366 -36092 386 -31858
rect -386 -36120 386 -36092
<< via3 >>
rect 302 31858 366 36092
rect 302 27328 366 31562
rect 302 22798 366 27032
rect 302 18268 366 22502
rect 302 13738 366 17972
rect 302 9208 366 13442
rect 302 4678 366 8912
rect 302 148 366 4382
rect 302 -4382 366 -148
rect 302 -8912 366 -4678
rect 302 -13442 366 -9208
rect 302 -17972 366 -13738
rect 302 -22502 366 -18268
rect 302 -27032 366 -22798
rect 302 -31562 366 -27328
rect 302 -36092 366 -31858
<< mimcap >>
rect -346 36040 54 36080
rect -346 31910 -306 36040
rect 14 31910 54 36040
rect -346 31870 54 31910
rect -346 31510 54 31550
rect -346 27380 -306 31510
rect 14 27380 54 31510
rect -346 27340 54 27380
rect -346 26980 54 27020
rect -346 22850 -306 26980
rect 14 22850 54 26980
rect -346 22810 54 22850
rect -346 22450 54 22490
rect -346 18320 -306 22450
rect 14 18320 54 22450
rect -346 18280 54 18320
rect -346 17920 54 17960
rect -346 13790 -306 17920
rect 14 13790 54 17920
rect -346 13750 54 13790
rect -346 13390 54 13430
rect -346 9260 -306 13390
rect 14 9260 54 13390
rect -346 9220 54 9260
rect -346 8860 54 8900
rect -346 4730 -306 8860
rect 14 4730 54 8860
rect -346 4690 54 4730
rect -346 4330 54 4370
rect -346 200 -306 4330
rect 14 200 54 4330
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -4330 -306 -200
rect 14 -4330 54 -200
rect -346 -4370 54 -4330
rect -346 -4730 54 -4690
rect -346 -8860 -306 -4730
rect 14 -8860 54 -4730
rect -346 -8900 54 -8860
rect -346 -9260 54 -9220
rect -346 -13390 -306 -9260
rect 14 -13390 54 -9260
rect -346 -13430 54 -13390
rect -346 -13790 54 -13750
rect -346 -17920 -306 -13790
rect 14 -17920 54 -13790
rect -346 -17960 54 -17920
rect -346 -18320 54 -18280
rect -346 -22450 -306 -18320
rect 14 -22450 54 -18320
rect -346 -22490 54 -22450
rect -346 -22850 54 -22810
rect -346 -26980 -306 -22850
rect 14 -26980 54 -22850
rect -346 -27020 54 -26980
rect -346 -27380 54 -27340
rect -346 -31510 -306 -27380
rect 14 -31510 54 -27380
rect -346 -31550 54 -31510
rect -346 -31910 54 -31870
rect -346 -36040 -306 -31910
rect 14 -36040 54 -31910
rect -346 -36080 54 -36040
<< mimcapcontact >>
rect -306 31910 14 36040
rect -306 27380 14 31510
rect -306 22850 14 26980
rect -306 18320 14 22450
rect -306 13790 14 17920
rect -306 9260 14 13390
rect -306 4730 14 8860
rect -306 200 14 4330
rect -306 -4330 14 -200
rect -306 -8860 14 -4730
rect -306 -13390 14 -9260
rect -306 -17920 14 -13790
rect -306 -22450 14 -18320
rect -306 -26980 14 -22850
rect -306 -31510 14 -27380
rect -306 -36040 14 -31910
<< metal4 >>
rect -198 36041 -94 36240
rect 282 36092 386 36240
rect -307 36040 15 36041
rect -307 31910 -306 36040
rect 14 31910 15 36040
rect -307 31909 15 31910
rect -198 31511 -94 31909
rect 282 31858 302 36092
rect 366 31858 386 36092
rect 282 31562 386 31858
rect -307 31510 15 31511
rect -307 27380 -306 31510
rect 14 27380 15 31510
rect -307 27379 15 27380
rect -198 26981 -94 27379
rect 282 27328 302 31562
rect 366 27328 386 31562
rect 282 27032 386 27328
rect -307 26980 15 26981
rect -307 22850 -306 26980
rect 14 22850 15 26980
rect -307 22849 15 22850
rect -198 22451 -94 22849
rect 282 22798 302 27032
rect 366 22798 386 27032
rect 282 22502 386 22798
rect -307 22450 15 22451
rect -307 18320 -306 22450
rect 14 18320 15 22450
rect -307 18319 15 18320
rect -198 17921 -94 18319
rect 282 18268 302 22502
rect 366 18268 386 22502
rect 282 17972 386 18268
rect -307 17920 15 17921
rect -307 13790 -306 17920
rect 14 13790 15 17920
rect -307 13789 15 13790
rect -198 13391 -94 13789
rect 282 13738 302 17972
rect 366 13738 386 17972
rect 282 13442 386 13738
rect -307 13390 15 13391
rect -307 9260 -306 13390
rect 14 9260 15 13390
rect -307 9259 15 9260
rect -198 8861 -94 9259
rect 282 9208 302 13442
rect 366 9208 386 13442
rect 282 8912 386 9208
rect -307 8860 15 8861
rect -307 4730 -306 8860
rect 14 4730 15 8860
rect -307 4729 15 4730
rect -198 4331 -94 4729
rect 282 4678 302 8912
rect 366 4678 386 8912
rect 282 4382 386 4678
rect -307 4330 15 4331
rect -307 200 -306 4330
rect 14 200 15 4330
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 4382
rect 366 148 386 4382
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -4330 -306 -200
rect 14 -4330 15 -200
rect -307 -4331 15 -4330
rect -198 -4729 -94 -4331
rect 282 -4382 302 -148
rect 366 -4382 386 -148
rect 282 -4678 386 -4382
rect -307 -4730 15 -4729
rect -307 -8860 -306 -4730
rect 14 -8860 15 -4730
rect -307 -8861 15 -8860
rect -198 -9259 -94 -8861
rect 282 -8912 302 -4678
rect 366 -8912 386 -4678
rect 282 -9208 386 -8912
rect -307 -9260 15 -9259
rect -307 -13390 -306 -9260
rect 14 -13390 15 -9260
rect -307 -13391 15 -13390
rect -198 -13789 -94 -13391
rect 282 -13442 302 -9208
rect 366 -13442 386 -9208
rect 282 -13738 386 -13442
rect -307 -13790 15 -13789
rect -307 -17920 -306 -13790
rect 14 -17920 15 -13790
rect -307 -17921 15 -17920
rect -198 -18319 -94 -17921
rect 282 -17972 302 -13738
rect 366 -17972 386 -13738
rect 282 -18268 386 -17972
rect -307 -18320 15 -18319
rect -307 -22450 -306 -18320
rect 14 -22450 15 -18320
rect -307 -22451 15 -22450
rect -198 -22849 -94 -22451
rect 282 -22502 302 -18268
rect 366 -22502 386 -18268
rect 282 -22798 386 -22502
rect -307 -22850 15 -22849
rect -307 -26980 -306 -22850
rect 14 -26980 15 -22850
rect -307 -26981 15 -26980
rect -198 -27379 -94 -26981
rect 282 -27032 302 -22798
rect 366 -27032 386 -22798
rect 282 -27328 386 -27032
rect -307 -27380 15 -27379
rect -307 -31510 -306 -27380
rect 14 -31510 15 -27380
rect -307 -31511 15 -31510
rect -198 -31909 -94 -31511
rect 282 -31562 302 -27328
rect 366 -31562 386 -27328
rect 282 -31858 386 -31562
rect -307 -31910 15 -31909
rect -307 -36040 -306 -31910
rect 14 -36040 15 -31910
rect -307 -36041 15 -36040
rect -198 -36240 -94 -36041
rect 282 -36092 302 -31858
rect 366 -36092 386 -31858
rect 282 -36240 386 -36092
<< properties >>
string FIXED_BBOX -386 31830 94 36120
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
