magic
tech sky130A
magscale 1 2
timestamp 1666052912
<< metal4 >>
rect -2047 2759 -949 2800
rect -2047 1081 -1205 2759
rect -969 1081 -949 2759
rect -2047 1040 -949 1081
rect -549 2759 549 2800
rect -549 1081 293 2759
rect 529 1081 549 2759
rect -549 1040 549 1081
rect 949 2759 2047 2800
rect 949 1081 1791 2759
rect 2027 1081 2047 2759
rect 949 1040 2047 1081
rect -2047 839 -949 880
rect -2047 -839 -1205 839
rect -969 -839 -949 839
rect -2047 -880 -949 -839
rect -549 839 549 880
rect -549 -839 293 839
rect 529 -839 549 839
rect -549 -880 549 -839
rect 949 839 2047 880
rect 949 -839 1791 839
rect 2027 -839 2047 839
rect 949 -880 2047 -839
rect -2047 -1081 -949 -1040
rect -2047 -2759 -1205 -1081
rect -969 -2759 -949 -1081
rect -2047 -2800 -949 -2759
rect -549 -1081 549 -1040
rect -549 -2759 293 -1081
rect 529 -2759 549 -1081
rect -549 -2800 549 -2759
rect 949 -1081 2047 -1040
rect 949 -2759 1791 -1081
rect 2027 -2759 2047 -1081
rect 949 -2800 2047 -2759
<< via4 >>
rect -1205 1081 -969 2759
rect 293 1081 529 2759
rect 1791 1081 2027 2759
rect -1205 -839 -969 839
rect 293 -839 529 839
rect 1791 -839 2027 839
rect -1205 -2759 -969 -1081
rect 293 -2759 529 -1081
rect 1791 -2759 2027 -1081
<< mimcap2 >>
rect -1967 2680 -1567 2720
rect -1967 1160 -1927 2680
rect -1607 1160 -1567 2680
rect -1967 1120 -1567 1160
rect -469 2680 -69 2720
rect -469 1160 -429 2680
rect -109 1160 -69 2680
rect -469 1120 -69 1160
rect 1029 2680 1429 2720
rect 1029 1160 1069 2680
rect 1389 1160 1429 2680
rect 1029 1120 1429 1160
rect -1967 760 -1567 800
rect -1967 -760 -1927 760
rect -1607 -760 -1567 760
rect -1967 -800 -1567 -760
rect -469 760 -69 800
rect -469 -760 -429 760
rect -109 -760 -69 760
rect -469 -800 -69 -760
rect 1029 760 1429 800
rect 1029 -760 1069 760
rect 1389 -760 1429 760
rect 1029 -800 1429 -760
rect -1967 -1160 -1567 -1120
rect -1967 -2680 -1927 -1160
rect -1607 -2680 -1567 -1160
rect -1967 -2720 -1567 -2680
rect -469 -1160 -69 -1120
rect -469 -2680 -429 -1160
rect -109 -2680 -69 -1160
rect -469 -2720 -69 -2680
rect 1029 -1160 1429 -1120
rect 1029 -2680 1069 -1160
rect 1389 -2680 1429 -1160
rect 1029 -2720 1429 -2680
<< mimcap2contact >>
rect -1927 1160 -1607 2680
rect -429 1160 -109 2680
rect 1069 1160 1389 2680
rect -1927 -760 -1607 760
rect -429 -760 -109 760
rect 1069 -760 1389 760
rect -1927 -2680 -1607 -1160
rect -429 -2680 -109 -1160
rect 1069 -2680 1389 -1160
<< metal5 >>
rect -1927 2704 -1607 2880
rect -1247 2759 -927 2880
rect -1951 2680 -1583 2704
rect -1951 1160 -1927 2680
rect -1607 1160 -1583 2680
rect -1951 1136 -1583 1160
rect -1927 784 -1607 1136
rect -1247 1081 -1205 2759
rect -969 1081 -927 2759
rect -429 2704 -109 2880
rect 251 2759 571 2880
rect -453 2680 -85 2704
rect -453 1160 -429 2680
rect -109 1160 -85 2680
rect -453 1136 -85 1160
rect -1247 839 -927 1081
rect -1951 760 -1583 784
rect -1951 -760 -1927 760
rect -1607 -760 -1583 760
rect -1951 -784 -1583 -760
rect -1927 -1136 -1607 -784
rect -1247 -839 -1205 839
rect -969 -839 -927 839
rect -429 784 -109 1136
rect 251 1081 293 2759
rect 529 1081 571 2759
rect 1069 2704 1389 2880
rect 1749 2759 2069 2880
rect 1045 2680 1413 2704
rect 1045 1160 1069 2680
rect 1389 1160 1413 2680
rect 1045 1136 1413 1160
rect 251 839 571 1081
rect -453 760 -85 784
rect -453 -760 -429 760
rect -109 -760 -85 760
rect -453 -784 -85 -760
rect -1247 -1081 -927 -839
rect -1951 -1160 -1583 -1136
rect -1951 -2680 -1927 -1160
rect -1607 -2680 -1583 -1160
rect -1951 -2704 -1583 -2680
rect -1927 -2880 -1607 -2704
rect -1247 -2759 -1205 -1081
rect -969 -2759 -927 -1081
rect -429 -1136 -109 -784
rect 251 -839 293 839
rect 529 -839 571 839
rect 1069 784 1389 1136
rect 1749 1081 1791 2759
rect 2027 1081 2069 2759
rect 1749 839 2069 1081
rect 1045 760 1413 784
rect 1045 -760 1069 760
rect 1389 -760 1413 760
rect 1045 -784 1413 -760
rect 251 -1081 571 -839
rect -453 -1160 -85 -1136
rect -453 -2680 -429 -1160
rect -109 -2680 -85 -1160
rect -453 -2704 -85 -2680
rect -1247 -2880 -927 -2759
rect -429 -2880 -109 -2704
rect 251 -2759 293 -1081
rect 529 -2759 571 -1081
rect 1069 -1136 1389 -784
rect 1749 -839 1791 839
rect 2027 -839 2069 839
rect 1749 -1081 2069 -839
rect 1045 -1160 1413 -1136
rect 1045 -2680 1069 -1160
rect 1389 -2680 1413 -1160
rect 1045 -2704 1413 -2680
rect 251 -2880 571 -2759
rect 1069 -2880 1389 -2704
rect 1749 -2759 1791 -1081
rect 2027 -2759 2069 -1081
rect 1749 -2880 2069 -2759
<< properties >>
string FIXED_BBOX 949 1040 1509 2800
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 2.00 l 8 val 35.8 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
