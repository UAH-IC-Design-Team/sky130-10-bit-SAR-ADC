magic
tech sky130A
magscale 1 2
timestamp 1666052912
<< metal3 >>
rect -948 792 -356 820
rect -948 368 -440 792
rect -376 368 -356 792
rect -948 340 -356 368
rect -296 792 296 820
rect -296 368 212 792
rect 276 368 296 792
rect -296 340 296 368
rect 356 792 948 820
rect 356 368 864 792
rect 928 368 948 792
rect 356 340 948 368
rect -948 212 -356 240
rect -948 -212 -440 212
rect -376 -212 -356 212
rect -948 -240 -356 -212
rect -296 212 296 240
rect -296 -212 212 212
rect 276 -212 296 212
rect -296 -240 296 -212
rect 356 212 948 240
rect 356 -212 864 212
rect 928 -212 948 212
rect 356 -240 948 -212
rect -948 -368 -356 -340
rect -948 -792 -440 -368
rect -376 -792 -356 -368
rect -948 -820 -356 -792
rect -296 -368 296 -340
rect -296 -792 212 -368
rect 276 -792 296 -368
rect -296 -820 296 -792
rect 356 -368 948 -340
rect 356 -792 864 -368
rect 928 -792 948 -368
rect 356 -820 948 -792
<< via3 >>
rect -440 368 -376 792
rect 212 368 276 792
rect 864 368 928 792
rect -440 -212 -376 212
rect 212 -212 276 212
rect 864 -212 928 212
rect -440 -792 -376 -368
rect 212 -792 276 -368
rect 864 -792 928 -368
<< mimcap >>
rect -908 740 -508 780
rect -908 420 -868 740
rect -548 420 -508 740
rect -908 380 -508 420
rect -256 740 144 780
rect -256 420 -216 740
rect 104 420 144 740
rect -256 380 144 420
rect 396 740 796 780
rect 396 420 436 740
rect 756 420 796 740
rect 396 380 796 420
rect -908 160 -508 200
rect -908 -160 -868 160
rect -548 -160 -508 160
rect -908 -200 -508 -160
rect -256 160 144 200
rect -256 -160 -216 160
rect 104 -160 144 160
rect -256 -200 144 -160
rect 396 160 796 200
rect 396 -160 436 160
rect 756 -160 796 160
rect 396 -200 796 -160
rect -908 -420 -508 -380
rect -908 -740 -868 -420
rect -548 -740 -508 -420
rect -908 -780 -508 -740
rect -256 -420 144 -380
rect -256 -740 -216 -420
rect 104 -740 144 -420
rect -256 -780 144 -740
rect 396 -420 796 -380
rect 396 -740 436 -420
rect 756 -740 796 -420
rect 396 -780 796 -740
<< mimcapcontact >>
rect -868 420 -548 740
rect -216 420 104 740
rect 436 420 756 740
rect -868 -160 -548 160
rect -216 -160 104 160
rect 436 -160 756 160
rect -868 -740 -548 -420
rect -216 -740 104 -420
rect 436 -740 756 -420
<< metal4 >>
rect -760 741 -656 870
rect -460 792 -356 870
rect -869 740 -547 741
rect -869 420 -868 740
rect -548 420 -547 740
rect -869 419 -547 420
rect -760 161 -656 419
rect -460 368 -440 792
rect -376 368 -356 792
rect -108 741 -4 870
rect 192 792 296 870
rect -217 740 105 741
rect -217 420 -216 740
rect 104 420 105 740
rect -217 419 105 420
rect -460 212 -356 368
rect -869 160 -547 161
rect -869 -160 -868 160
rect -548 -160 -547 160
rect -869 -161 -547 -160
rect -760 -419 -656 -161
rect -460 -212 -440 212
rect -376 -212 -356 212
rect -108 161 -4 419
rect 192 368 212 792
rect 276 368 296 792
rect 544 741 648 870
rect 844 792 948 870
rect 435 740 757 741
rect 435 420 436 740
rect 756 420 757 740
rect 435 419 757 420
rect 192 212 296 368
rect -217 160 105 161
rect -217 -160 -216 160
rect 104 -160 105 160
rect -217 -161 105 -160
rect -460 -368 -356 -212
rect -869 -420 -547 -419
rect -869 -740 -868 -420
rect -548 -740 -547 -420
rect -869 -741 -547 -740
rect -760 -870 -656 -741
rect -460 -792 -440 -368
rect -376 -792 -356 -368
rect -108 -419 -4 -161
rect 192 -212 212 212
rect 276 -212 296 212
rect 544 161 648 419
rect 844 368 864 792
rect 928 368 948 792
rect 844 212 948 368
rect 435 160 757 161
rect 435 -160 436 160
rect 756 -160 757 160
rect 435 -161 757 -160
rect 192 -368 296 -212
rect -217 -420 105 -419
rect -217 -740 -216 -420
rect 104 -740 105 -420
rect -217 -741 105 -740
rect -460 -870 -356 -792
rect -108 -870 -4 -741
rect 192 -792 212 -368
rect 276 -792 296 -368
rect 544 -419 648 -161
rect 844 -212 864 212
rect 928 -212 948 212
rect 844 -368 948 -212
rect 435 -420 757 -419
rect 435 -740 436 -420
rect 756 -740 757 -420
rect 435 -741 757 -740
rect 192 -870 296 -792
rect 544 -870 648 -741
rect 844 -792 864 -368
rect 928 -792 948 -368
rect 844 -870 948 -792
<< properties >>
string FIXED_BBOX 356 340 836 820
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
