magic
tech sky130A
magscale 1 2
timestamp 1667436771
<< error_p >>
rect -119 62 -73 74
rect 73 62 119 74
rect -119 28 -113 62
rect 73 28 79 62
rect -119 16 -73 28
rect 73 16 119 28
rect -215 -28 -169 -16
rect -23 -28 23 -16
rect 169 -28 215 -16
rect -215 -62 -209 -28
rect -23 -62 -17 -28
rect 169 -62 175 -28
rect -215 -74 -169 -62
rect -23 -74 23 -62
rect 169 -74 215 -62
<< nmos >>
rect -159 -91 -129 91
rect -63 -91 -33 91
rect 33 -91 63 91
rect 129 -91 159 91
<< ndiff >>
rect -221 79 -159 91
rect -221 -79 -209 79
rect -175 -79 -159 79
rect -221 -91 -159 -79
rect -129 79 -63 91
rect -129 -79 -113 79
rect -79 -79 -63 79
rect -129 -91 -63 -79
rect -33 79 33 91
rect -33 -79 -17 79
rect 17 -79 33 79
rect -33 -91 33 -79
rect 63 79 129 91
rect 63 -79 79 79
rect 113 -79 129 79
rect 63 -91 129 -79
rect 159 79 221 91
rect 159 -79 175 79
rect 209 -79 221 79
rect 159 -91 221 -79
<< ndiffc >>
rect -209 -79 -175 79
rect -113 -79 -79 79
rect -17 -79 17 79
rect 79 -79 113 79
rect 175 -79 209 79
<< poly >>
rect -159 91 -129 119
rect -63 91 -33 119
rect 33 91 63 119
rect 129 91 159 119
rect -159 -113 -129 -91
rect -63 -113 -33 -91
rect 33 -113 63 -91
rect 129 -113 159 -91
rect -177 -129 189 -113
rect -177 -163 -161 -129
rect -127 -163 -66 -129
rect -32 -163 31 -129
rect 65 -163 124 -129
rect 158 -163 189 -129
rect -177 -179 189 -163
<< polycont >>
rect -161 -163 -127 -129
rect -66 -163 -32 -129
rect 31 -163 65 -129
rect 124 -163 158 -129
<< locali >>
rect -209 79 -175 95
rect -209 -95 -175 -79
rect -113 79 -79 95
rect -113 -95 -79 -79
rect -17 79 17 95
rect -17 -95 17 -79
rect 79 79 113 95
rect 79 -95 113 -79
rect 175 79 209 95
rect 175 -95 209 -79
rect -177 -163 -161 -129
rect -127 -163 -66 -129
rect -32 -163 31 -129
rect 65 -163 124 -129
rect 158 -163 189 -129
<< viali >>
rect -209 -62 -175 -28
rect -113 28 -79 62
rect -17 -62 17 -28
rect 79 28 113 62
rect 175 -62 209 -28
rect -161 -163 -127 -129
rect -66 -163 -32 -129
rect 31 -163 65 -129
rect 124 -163 158 -129
<< metal1 >>
rect -119 62 -73 74
rect -119 28 -113 62
rect -79 28 -73 62
rect -119 16 -73 28
rect 73 62 119 74
rect 73 28 79 62
rect 113 28 119 62
rect 73 16 119 28
rect -215 -28 -169 -16
rect -215 -62 -209 -28
rect -175 -62 -169 -28
rect -215 -74 -169 -62
rect -23 -28 23 -16
rect -23 -62 -17 -28
rect 17 -62 23 -28
rect -23 -74 23 -62
rect 169 -28 215 -16
rect 169 -62 175 -28
rect 209 -62 215 -28
rect 169 -74 215 -62
rect -177 -129 189 -123
rect -177 -163 -161 -129
rect -127 -163 -66 -129
rect -32 -163 31 -129
rect 65 -163 124 -129
rect 158 -163 189 -129
rect -177 -169 189 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc -20 viadrn +20 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
