magic
tech sky130A
timestamp 1667684479
<< metal4 >>
rect 250 5200 310 5800
rect 590 5200 650 5800
rect 250 4400 310 5000
rect 590 4400 650 5000
rect 250 3600 310 4200
rect 590 3600 650 4200
rect 250 2800 310 3400
rect 590 2800 650 3400
rect 250 2000 310 2600
rect 590 2000 650 2600
rect 250 1200 310 1800
rect 590 1200 650 1800
rect 250 400 310 1000
rect 590 400 650 1000
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
array 0 0 800 0 7 800
timestamp 1667663783
transform 1 0 325 0 1 300
box -325 -300 325 300
<< end >>
