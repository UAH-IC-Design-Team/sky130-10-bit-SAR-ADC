magic
tech sky130A
magscale 1 2
timestamp 1667868455
<< pwell >>
rect 420 20 600 210
<< ndiode >>
rect 447 167 573 185
rect 447 133 456 167
rect 490 133 531 167
rect 565 133 573 167
rect 447 99 573 133
rect 447 65 456 99
rect 490 65 531 99
rect 565 65 573 99
rect 447 47 573 65
<< ndiodec >>
rect 456 133 490 167
rect 531 133 565 167
rect 456 65 490 99
rect 531 65 565 99
<< locali >>
rect 430 190 590 200
rect 430 40 440 190
rect 580 40 590 190
rect 430 30 590 40
<< viali >>
rect 440 167 580 190
rect 440 133 456 167
rect 456 133 490 167
rect 490 133 531 167
rect 531 133 565 167
rect 565 133 580 167
rect 440 99 580 133
rect 440 65 456 99
rect 456 65 490 99
rect 490 65 531 99
rect 531 65 565 99
rect 565 65 580 99
rect 440 40 580 65
<< metal1 >>
rect 420 190 600 210
rect 420 40 440 190
rect 580 40 600 190
rect 420 20 600 40
<< end >>
