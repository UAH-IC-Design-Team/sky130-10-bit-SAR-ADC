* NGSPICE file created from demux2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_0 A B VGND VPWR X VNB VPB a_40_47#
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.795e+11p pd=3.89e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.696e+11p pd=1.81e+06u as=0p ps=0u w=640000u l=150000u
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=1.932e+11p pd=1.76e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=150000u
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt demux2 VDD VSS S IN OUT_0 OUT_1
Xx1 x3/Y IN VSS VDD OUT_0 VSS VDD x1/a_40_47# sky130_fd_sc_hd__and2_0
Xx2 S IN VSS VDD OUT_1 VSS VDD x2/a_40_47# sky130_fd_sc_hd__and2_0
Xx3 S VSS VDD x3/Y VSS VDD sky130_fd_sc_hd__inv_1
.ends

