magic
tech sky130A
magscale 1 2
timestamp 1667435063
<< nmos >>
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
<< ndiff >>
rect -509 488 -447 500
rect -509 -488 -497 488
rect -463 -488 -447 488
rect -509 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 509 500
rect 447 -488 463 488
rect 497 -488 509 488
rect 447 -500 509 -488
<< ndiffc >>
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
<< poly >>
rect -465 582 481 598
rect -465 548 -449 582
rect -415 548 -354 582
rect -320 548 -257 582
rect -223 548 -164 582
rect -130 548 -65 582
rect -31 548 26 582
rect 60 548 127 582
rect 161 548 216 582
rect 250 548 319 582
rect 353 548 416 582
rect 450 548 481 582
rect -465 532 481 548
rect -447 500 -417 532
rect -351 500 -321 532
rect -255 500 -225 532
rect -159 500 -129 532
rect -63 500 -33 532
rect 33 500 63 532
rect 129 500 159 532
rect 225 500 255 532
rect 321 500 351 532
rect 417 500 447 532
rect -447 -532 -417 -500
rect -351 -532 -321 -500
rect -255 -532 -225 -500
rect -159 -532 -129 -500
rect -63 -532 -33 -500
rect 33 -532 63 -500
rect 129 -532 159 -500
rect 225 -532 255 -500
rect 321 -532 351 -500
rect 417 -532 447 -500
<< polycont >>
rect -449 548 -415 582
rect -354 548 -320 582
rect -257 548 -223 582
rect -164 548 -130 582
rect -65 548 -31 582
rect 26 548 60 582
rect 127 548 161 582
rect 216 548 250 582
rect 319 548 353 582
rect 416 548 450 582
<< locali >>
rect -465 548 -449 582
rect -415 548 -354 582
rect -320 548 -257 582
rect -223 548 -164 582
rect -130 548 -65 582
rect -31 548 26 582
rect 60 548 127 582
rect 161 548 216 582
rect 250 548 319 582
rect 353 548 416 582
rect 450 548 481 582
rect -497 488 -463 504
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect 463 488 497 504
rect 463 -504 497 -488
<< viali >>
rect -449 548 -415 582
rect -354 548 -320 582
rect -257 548 -223 582
rect -164 548 -130 582
rect -65 548 -31 582
rect 26 548 60 582
rect 127 548 161 582
rect 216 548 250 582
rect 319 548 353 582
rect 416 548 450 582
rect -497 -471 -463 -81
rect -401 81 -367 471
rect -305 -471 -271 -81
rect -209 81 -175 471
rect -113 -471 -79 -81
rect -17 81 17 471
rect 79 -471 113 -81
rect 175 81 209 471
rect 271 -471 305 -81
rect 367 81 401 471
rect 463 -471 497 -81
<< metal1 >>
rect -465 582 481 588
rect -465 548 -449 582
rect -415 548 -354 582
rect -320 548 -257 582
rect -223 548 -164 582
rect -130 548 -65 582
rect -31 548 26 582
rect 60 548 127 582
rect 161 548 216 582
rect 250 548 319 582
rect 353 548 416 582
rect 450 548 481 582
rect -465 542 481 548
rect -407 471 -361 483
rect -407 81 -401 471
rect -367 81 -361 471
rect -407 69 -361 81
rect -215 471 -169 483
rect -215 81 -209 471
rect -175 81 -169 471
rect -215 69 -169 81
rect -23 471 23 483
rect -23 81 -17 471
rect 17 81 23 471
rect -23 69 23 81
rect 169 471 215 483
rect 169 81 175 471
rect 209 81 215 471
rect 169 69 215 81
rect 361 471 407 483
rect 361 81 367 471
rect 401 81 407 471
rect 361 69 407 81
rect -503 -81 -457 -69
rect -503 -471 -497 -81
rect -463 -471 -457 -81
rect -503 -483 -457 -471
rect -311 -81 -265 -69
rect -311 -471 -305 -81
rect -271 -471 -265 -81
rect -311 -483 -265 -471
rect -119 -81 -73 -69
rect -119 -471 -113 -81
rect -79 -471 -73 -81
rect -119 -483 -73 -471
rect 73 -81 119 -69
rect 73 -471 79 -81
rect 113 -471 119 -81
rect 73 -483 119 -471
rect 265 -81 311 -69
rect 265 -471 271 -81
rect 305 -471 311 -81
rect 265 -483 311 -471
rect 457 -81 503 -69
rect 457 -471 463 -81
rect 497 -471 503 -81
rect 457 -483 503 -471
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
