magic
tech sky130A
magscale 1 2
timestamp 1666649035
<< error_p >>
rect -605 527 -547 533
rect -413 527 -355 533
rect -221 527 -163 533
rect -29 527 29 533
rect 163 527 221 533
rect 355 527 413 533
rect 547 527 605 533
rect -605 493 -593 527
rect -413 493 -401 527
rect -221 493 -209 527
rect -29 493 -17 527
rect 163 493 175 527
rect 355 493 367 527
rect 547 493 559 527
rect -605 487 -547 493
rect -413 487 -355 493
rect -221 487 -163 493
rect -29 487 29 493
rect 163 487 221 493
rect 355 487 413 493
rect 547 487 605 493
rect -701 -493 -643 -487
rect -509 -493 -451 -487
rect -317 -493 -259 -487
rect -125 -493 -67 -487
rect 67 -493 125 -487
rect 259 -493 317 -487
rect 451 -493 509 -487
rect 643 -493 701 -487
rect -701 -527 -689 -493
rect -509 -527 -497 -493
rect -317 -527 -305 -493
rect -125 -527 -113 -493
rect 67 -527 79 -493
rect 259 -527 271 -493
rect 451 -527 463 -493
rect 643 -527 655 -493
rect -701 -533 -643 -527
rect -509 -533 -451 -527
rect -317 -533 -259 -527
rect -125 -533 -67 -527
rect 67 -533 125 -527
rect 259 -533 317 -527
rect 451 -533 509 -527
rect 643 -533 701 -527
<< pwell >>
rect -887 -665 887 665
<< nmos >>
rect -687 -455 -657 455
rect -591 -455 -561 455
rect -495 -455 -465 455
rect -399 -455 -369 455
rect -303 -455 -273 455
rect -207 -455 -177 455
rect -111 -455 -81 455
rect -15 -455 15 455
rect 81 -455 111 455
rect 177 -455 207 455
rect 273 -455 303 455
rect 369 -455 399 455
rect 465 -455 495 455
rect 561 -455 591 455
rect 657 -455 687 455
<< ndiff >>
rect -749 443 -687 455
rect -749 -443 -737 443
rect -703 -443 -687 443
rect -749 -455 -687 -443
rect -657 443 -591 455
rect -657 -443 -641 443
rect -607 -443 -591 443
rect -657 -455 -591 -443
rect -561 443 -495 455
rect -561 -443 -545 443
rect -511 -443 -495 443
rect -561 -455 -495 -443
rect -465 443 -399 455
rect -465 -443 -449 443
rect -415 -443 -399 443
rect -465 -455 -399 -443
rect -369 443 -303 455
rect -369 -443 -353 443
rect -319 -443 -303 443
rect -369 -455 -303 -443
rect -273 443 -207 455
rect -273 -443 -257 443
rect -223 -443 -207 443
rect -273 -455 -207 -443
rect -177 443 -111 455
rect -177 -443 -161 443
rect -127 -443 -111 443
rect -177 -455 -111 -443
rect -81 443 -15 455
rect -81 -443 -65 443
rect -31 -443 -15 443
rect -81 -455 -15 -443
rect 15 443 81 455
rect 15 -443 31 443
rect 65 -443 81 443
rect 15 -455 81 -443
rect 111 443 177 455
rect 111 -443 127 443
rect 161 -443 177 443
rect 111 -455 177 -443
rect 207 443 273 455
rect 207 -443 223 443
rect 257 -443 273 443
rect 207 -455 273 -443
rect 303 443 369 455
rect 303 -443 319 443
rect 353 -443 369 443
rect 303 -455 369 -443
rect 399 443 465 455
rect 399 -443 415 443
rect 449 -443 465 443
rect 399 -455 465 -443
rect 495 443 561 455
rect 495 -443 511 443
rect 545 -443 561 443
rect 495 -455 561 -443
rect 591 443 657 455
rect 591 -443 607 443
rect 641 -443 657 443
rect 591 -455 657 -443
rect 687 443 749 455
rect 687 -443 703 443
rect 737 -443 749 443
rect 687 -455 749 -443
<< ndiffc >>
rect -737 -443 -703 443
rect -641 -443 -607 443
rect -545 -443 -511 443
rect -449 -443 -415 443
rect -353 -443 -319 443
rect -257 -443 -223 443
rect -161 -443 -127 443
rect -65 -443 -31 443
rect 31 -443 65 443
rect 127 -443 161 443
rect 223 -443 257 443
rect 319 -443 353 443
rect 415 -443 449 443
rect 511 -443 545 443
rect 607 -443 641 443
rect 703 -443 737 443
<< psubdiff >>
rect -851 595 -755 629
rect 755 595 851 629
rect -851 533 -817 595
rect 817 533 851 595
rect -851 -595 -817 -533
rect 817 -595 851 -533
rect -851 -629 -755 -595
rect 755 -629 851 -595
<< psubdiffcont >>
rect -755 595 755 629
rect -851 -533 -817 533
rect 817 -533 851 533
rect -755 -629 755 -595
<< poly >>
rect -609 527 -543 543
rect -609 493 -593 527
rect -559 493 -543 527
rect -687 455 -657 481
rect -609 477 -543 493
rect -417 527 -351 543
rect -417 493 -401 527
rect -367 493 -351 527
rect -591 455 -561 477
rect -495 455 -465 481
rect -417 477 -351 493
rect -225 527 -159 543
rect -225 493 -209 527
rect -175 493 -159 527
rect -399 455 -369 477
rect -303 455 -273 481
rect -225 477 -159 493
rect -33 527 33 543
rect -33 493 -17 527
rect 17 493 33 527
rect -207 455 -177 477
rect -111 455 -81 481
rect -33 477 33 493
rect 159 527 225 543
rect 159 493 175 527
rect 209 493 225 527
rect -15 455 15 477
rect 81 455 111 481
rect 159 477 225 493
rect 351 527 417 543
rect 351 493 367 527
rect 401 493 417 527
rect 177 455 207 477
rect 273 455 303 481
rect 351 477 417 493
rect 543 527 609 543
rect 543 493 559 527
rect 593 493 609 527
rect 369 455 399 477
rect 465 455 495 481
rect 543 477 609 493
rect 561 455 591 477
rect 657 455 687 481
rect -687 -477 -657 -455
rect -705 -493 -639 -477
rect -591 -481 -561 -455
rect -495 -477 -465 -455
rect -705 -527 -689 -493
rect -655 -527 -639 -493
rect -705 -543 -639 -527
rect -513 -493 -447 -477
rect -399 -481 -369 -455
rect -303 -477 -273 -455
rect -513 -527 -497 -493
rect -463 -527 -447 -493
rect -513 -543 -447 -527
rect -321 -493 -255 -477
rect -207 -481 -177 -455
rect -111 -477 -81 -455
rect -321 -527 -305 -493
rect -271 -527 -255 -493
rect -321 -543 -255 -527
rect -129 -493 -63 -477
rect -15 -481 15 -455
rect 81 -477 111 -455
rect -129 -527 -113 -493
rect -79 -527 -63 -493
rect -129 -543 -63 -527
rect 63 -493 129 -477
rect 177 -481 207 -455
rect 273 -477 303 -455
rect 63 -527 79 -493
rect 113 -527 129 -493
rect 63 -543 129 -527
rect 255 -493 321 -477
rect 369 -481 399 -455
rect 465 -477 495 -455
rect 255 -527 271 -493
rect 305 -527 321 -493
rect 255 -543 321 -527
rect 447 -493 513 -477
rect 561 -481 591 -455
rect 657 -477 687 -455
rect 447 -527 463 -493
rect 497 -527 513 -493
rect 447 -543 513 -527
rect 639 -493 705 -477
rect 639 -527 655 -493
rect 689 -527 705 -493
rect 639 -543 705 -527
<< polycont >>
rect -593 493 -559 527
rect -401 493 -367 527
rect -209 493 -175 527
rect -17 493 17 527
rect 175 493 209 527
rect 367 493 401 527
rect 559 493 593 527
rect -689 -527 -655 -493
rect -497 -527 -463 -493
rect -305 -527 -271 -493
rect -113 -527 -79 -493
rect 79 -527 113 -493
rect 271 -527 305 -493
rect 463 -527 497 -493
rect 655 -527 689 -493
<< locali >>
rect -851 595 -755 629
rect 755 595 851 629
rect -851 533 -817 595
rect 817 533 851 595
rect -609 493 -593 527
rect -559 493 -543 527
rect -417 493 -401 527
rect -367 493 -351 527
rect -225 493 -209 527
rect -175 493 -159 527
rect -33 493 -17 527
rect 17 493 33 527
rect 159 493 175 527
rect 209 493 225 527
rect 351 493 367 527
rect 401 493 417 527
rect 543 493 559 527
rect 593 493 609 527
rect -737 443 -703 459
rect -737 -459 -703 -443
rect -641 443 -607 459
rect -641 -459 -607 -443
rect -545 443 -511 459
rect -545 -459 -511 -443
rect -449 443 -415 459
rect -449 -459 -415 -443
rect -353 443 -319 459
rect -353 -459 -319 -443
rect -257 443 -223 459
rect -257 -459 -223 -443
rect -161 443 -127 459
rect -161 -459 -127 -443
rect -65 443 -31 459
rect -65 -459 -31 -443
rect 31 443 65 459
rect 31 -459 65 -443
rect 127 443 161 459
rect 127 -459 161 -443
rect 223 443 257 459
rect 223 -459 257 -443
rect 319 443 353 459
rect 319 -459 353 -443
rect 415 443 449 459
rect 415 -459 449 -443
rect 511 443 545 459
rect 511 -459 545 -443
rect 607 443 641 459
rect 607 -459 641 -443
rect 703 443 737 459
rect 703 -459 737 -443
rect -705 -527 -689 -493
rect -655 -527 -639 -493
rect -513 -527 -497 -493
rect -463 -527 -447 -493
rect -321 -527 -305 -493
rect -271 -527 -255 -493
rect -129 -527 -113 -493
rect -79 -527 -63 -493
rect 63 -527 79 -493
rect 113 -527 129 -493
rect 255 -527 271 -493
rect 305 -527 321 -493
rect 447 -527 463 -493
rect 497 -527 513 -493
rect 639 -527 655 -493
rect 689 -527 705 -493
rect -851 -595 -817 -533
rect 817 -595 851 -533
rect -851 -629 -755 -595
rect 755 -629 851 -595
<< viali >>
rect -593 493 -559 527
rect -401 493 -367 527
rect -209 493 -175 527
rect -17 493 17 527
rect 175 493 209 527
rect 367 493 401 527
rect 559 493 593 527
rect -737 -443 -703 443
rect -641 -443 -607 443
rect -545 -443 -511 443
rect -449 -443 -415 443
rect -353 -443 -319 443
rect -257 -443 -223 443
rect -161 -443 -127 443
rect -65 -443 -31 443
rect 31 -443 65 443
rect 127 -443 161 443
rect 223 -443 257 443
rect 319 -443 353 443
rect 415 -443 449 443
rect 511 -443 545 443
rect 607 -443 641 443
rect 703 -443 737 443
rect -689 -527 -655 -493
rect -497 -527 -463 -493
rect -305 -527 -271 -493
rect -113 -527 -79 -493
rect 79 -527 113 -493
rect 271 -527 305 -493
rect 463 -527 497 -493
rect 655 -527 689 -493
<< metal1 >>
rect -605 527 -547 533
rect -605 493 -593 527
rect -559 493 -547 527
rect -605 487 -547 493
rect -413 527 -355 533
rect -413 493 -401 527
rect -367 493 -355 527
rect -413 487 -355 493
rect -221 527 -163 533
rect -221 493 -209 527
rect -175 493 -163 527
rect -221 487 -163 493
rect -29 527 29 533
rect -29 493 -17 527
rect 17 493 29 527
rect -29 487 29 493
rect 163 527 221 533
rect 163 493 175 527
rect 209 493 221 527
rect 163 487 221 493
rect 355 527 413 533
rect 355 493 367 527
rect 401 493 413 527
rect 355 487 413 493
rect 547 527 605 533
rect 547 493 559 527
rect 593 493 605 527
rect 547 487 605 493
rect -743 443 -697 455
rect -743 -443 -737 443
rect -703 -443 -697 443
rect -743 -455 -697 -443
rect -647 443 -601 455
rect -647 -443 -641 443
rect -607 -443 -601 443
rect -647 -455 -601 -443
rect -551 443 -505 455
rect -551 -443 -545 443
rect -511 -443 -505 443
rect -551 -455 -505 -443
rect -455 443 -409 455
rect -455 -443 -449 443
rect -415 -443 -409 443
rect -455 -455 -409 -443
rect -359 443 -313 455
rect -359 -443 -353 443
rect -319 -443 -313 443
rect -359 -455 -313 -443
rect -263 443 -217 455
rect -263 -443 -257 443
rect -223 -443 -217 443
rect -263 -455 -217 -443
rect -167 443 -121 455
rect -167 -443 -161 443
rect -127 -443 -121 443
rect -167 -455 -121 -443
rect -71 443 -25 455
rect -71 -443 -65 443
rect -31 -443 -25 443
rect -71 -455 -25 -443
rect 25 443 71 455
rect 25 -443 31 443
rect 65 -443 71 443
rect 25 -455 71 -443
rect 121 443 167 455
rect 121 -443 127 443
rect 161 -443 167 443
rect 121 -455 167 -443
rect 217 443 263 455
rect 217 -443 223 443
rect 257 -443 263 443
rect 217 -455 263 -443
rect 313 443 359 455
rect 313 -443 319 443
rect 353 -443 359 443
rect 313 -455 359 -443
rect 409 443 455 455
rect 409 -443 415 443
rect 449 -443 455 443
rect 409 -455 455 -443
rect 505 443 551 455
rect 505 -443 511 443
rect 545 -443 551 443
rect 505 -455 551 -443
rect 601 443 647 455
rect 601 -443 607 443
rect 641 -443 647 443
rect 601 -455 647 -443
rect 697 443 743 455
rect 697 -443 703 443
rect 737 -443 743 443
rect 697 -455 743 -443
rect -701 -493 -643 -487
rect -701 -527 -689 -493
rect -655 -527 -643 -493
rect -701 -533 -643 -527
rect -509 -493 -451 -487
rect -509 -527 -497 -493
rect -463 -527 -451 -493
rect -509 -533 -451 -527
rect -317 -493 -259 -487
rect -317 -527 -305 -493
rect -271 -527 -259 -493
rect -317 -533 -259 -527
rect -125 -493 -67 -487
rect -125 -527 -113 -493
rect -79 -527 -67 -493
rect -125 -533 -67 -527
rect 67 -493 125 -487
rect 67 -527 79 -493
rect 113 -527 125 -493
rect 67 -533 125 -527
rect 259 -493 317 -487
rect 259 -527 271 -493
rect 305 -527 317 -493
rect 259 -533 317 -527
rect 451 -493 509 -487
rect 451 -527 463 -493
rect 497 -527 509 -493
rect 451 -533 509 -527
rect 643 -493 701 -487
rect 643 -527 655 -493
rect 689 -527 701 -493
rect 643 -533 701 -527
<< properties >>
string FIXED_BBOX -834 -612 834 612
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.55 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
