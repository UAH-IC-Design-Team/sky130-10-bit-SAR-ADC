magic
tech sky130A
magscale 1 2
timestamp 1666486738
<< error_p >>
rect -29 363 29 369
rect -29 329 -17 363
rect -29 323 29 329
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -329 29 -323
rect -29 -363 -17 -329
rect -29 -369 29 -363
<< nmos >>
rect -15 109 15 291
rect -15 -291 15 -109
<< ndiff >>
rect -73 279 -15 291
rect -73 121 -61 279
rect -27 121 -15 279
rect -73 109 -15 121
rect 15 279 73 291
rect 15 121 27 279
rect 61 121 73 279
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -279 -61 -121
rect -27 -279 -15 -121
rect -73 -291 -15 -279
rect 15 -121 73 -109
rect 15 -279 27 -121
rect 61 -279 73 -121
rect 15 -291 73 -279
<< ndiffc >>
rect -61 121 -27 279
rect 27 121 61 279
rect -61 -279 -27 -121
rect 27 -279 61 -121
<< poly >>
rect -33 363 33 379
rect -33 329 -17 363
rect 17 329 33 363
rect -33 313 33 329
rect -15 291 15 313
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -313 15 -291
rect -33 -329 33 -313
rect -33 -363 -17 -329
rect 17 -363 33 -329
rect -33 -379 33 -363
<< polycont >>
rect -17 329 17 363
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -363 17 -329
<< locali >>
rect -33 329 -17 363
rect 17 329 33 363
rect -61 279 -27 295
rect -61 105 -27 121
rect 27 279 61 295
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -295 -27 -279
rect 27 -121 61 -105
rect 27 -295 61 -279
rect -33 -363 -17 -329
rect 17 -363 33 -329
<< viali >>
rect -17 329 17 363
rect -61 121 -27 279
rect 27 121 61 279
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -279 -27 -121
rect 27 -279 61 -121
rect -17 -363 17 -329
<< metal1 >>
rect -29 363 29 369
rect -29 329 -17 363
rect 17 329 29 363
rect -29 323 29 329
rect -67 279 -21 291
rect -67 121 -61 279
rect -27 121 -21 279
rect -67 109 -21 121
rect 21 279 67 291
rect 21 121 27 279
rect 61 121 67 279
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -279 -61 -121
rect -27 -279 -21 -121
rect -67 -291 -21 -279
rect 21 -121 67 -109
rect 21 -279 27 -121
rect 61 -279 67 -121
rect 21 -291 67 -279
rect -29 -329 29 -323
rect -29 -363 -17 -329
rect 17 -363 29 -329
rect -29 -369 29 -363
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
