magic
tech sky130A
magscale 1 2
timestamp 1666552007
<< error_p >>
rect -29 1563 29 1569
rect -29 1529 -17 1563
rect -29 1523 29 1529
rect -29 1271 29 1277
rect -29 1237 -17 1271
rect -29 1231 29 1237
rect -29 1163 29 1169
rect -29 1129 -17 1163
rect -29 1123 29 1129
rect -29 871 29 877
rect -29 837 -17 871
rect -29 831 29 837
rect -29 763 29 769
rect -29 729 -17 763
rect -29 723 29 729
rect -29 471 29 477
rect -29 437 -17 471
rect -29 431 29 437
rect -29 363 29 369
rect -29 329 -17 363
rect -29 323 29 329
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -329 29 -323
rect -29 -363 -17 -329
rect -29 -369 29 -363
rect -29 -437 29 -431
rect -29 -471 -17 -437
rect -29 -477 29 -471
rect -29 -729 29 -723
rect -29 -763 -17 -729
rect -29 -769 29 -763
rect -29 -837 29 -831
rect -29 -871 -17 -837
rect -29 -877 29 -871
rect -29 -1129 29 -1123
rect -29 -1163 -17 -1129
rect -29 -1169 29 -1163
rect -29 -1237 29 -1231
rect -29 -1271 -17 -1237
rect -29 -1277 29 -1271
rect -29 -1529 29 -1523
rect -29 -1563 -17 -1529
rect -29 -1569 29 -1563
<< nmos >>
rect -15 1309 15 1491
rect -15 909 15 1091
rect -15 509 15 691
rect -15 109 15 291
rect -15 -291 15 -109
rect -15 -691 15 -509
rect -15 -1091 15 -909
rect -15 -1491 15 -1309
<< ndiff >>
rect -73 1479 -15 1491
rect -73 1321 -61 1479
rect -27 1321 -15 1479
rect -73 1309 -15 1321
rect 15 1479 73 1491
rect 15 1321 27 1479
rect 61 1321 73 1479
rect 15 1309 73 1321
rect -73 1079 -15 1091
rect -73 921 -61 1079
rect -27 921 -15 1079
rect -73 909 -15 921
rect 15 1079 73 1091
rect 15 921 27 1079
rect 61 921 73 1079
rect 15 909 73 921
rect -73 679 -15 691
rect -73 521 -61 679
rect -27 521 -15 679
rect -73 509 -15 521
rect 15 679 73 691
rect 15 521 27 679
rect 61 521 73 679
rect 15 509 73 521
rect -73 279 -15 291
rect -73 121 -61 279
rect -27 121 -15 279
rect -73 109 -15 121
rect 15 279 73 291
rect 15 121 27 279
rect 61 121 73 279
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -279 -61 -121
rect -27 -279 -15 -121
rect -73 -291 -15 -279
rect 15 -121 73 -109
rect 15 -279 27 -121
rect 61 -279 73 -121
rect 15 -291 73 -279
rect -73 -521 -15 -509
rect -73 -679 -61 -521
rect -27 -679 -15 -521
rect -73 -691 -15 -679
rect 15 -521 73 -509
rect 15 -679 27 -521
rect 61 -679 73 -521
rect 15 -691 73 -679
rect -73 -921 -15 -909
rect -73 -1079 -61 -921
rect -27 -1079 -15 -921
rect -73 -1091 -15 -1079
rect 15 -921 73 -909
rect 15 -1079 27 -921
rect 61 -1079 73 -921
rect 15 -1091 73 -1079
rect -73 -1321 -15 -1309
rect -73 -1479 -61 -1321
rect -27 -1479 -15 -1321
rect -73 -1491 -15 -1479
rect 15 -1321 73 -1309
rect 15 -1479 27 -1321
rect 61 -1479 73 -1321
rect 15 -1491 73 -1479
<< ndiffc >>
rect -61 1321 -27 1479
rect 27 1321 61 1479
rect -61 921 -27 1079
rect 27 921 61 1079
rect -61 521 -27 679
rect 27 521 61 679
rect -61 121 -27 279
rect 27 121 61 279
rect -61 -279 -27 -121
rect 27 -279 61 -121
rect -61 -679 -27 -521
rect 27 -679 61 -521
rect -61 -1079 -27 -921
rect 27 -1079 61 -921
rect -61 -1479 -27 -1321
rect 27 -1479 61 -1321
<< poly >>
rect -33 1563 33 1579
rect -33 1529 -17 1563
rect 17 1529 33 1563
rect -33 1513 33 1529
rect -15 1491 15 1513
rect -15 1287 15 1309
rect -33 1271 33 1287
rect -33 1237 -17 1271
rect 17 1237 33 1271
rect -33 1221 33 1237
rect -33 1163 33 1179
rect -33 1129 -17 1163
rect 17 1129 33 1163
rect -33 1113 33 1129
rect -15 1091 15 1113
rect -15 887 15 909
rect -33 871 33 887
rect -33 837 -17 871
rect 17 837 33 871
rect -33 821 33 837
rect -33 763 33 779
rect -33 729 -17 763
rect 17 729 33 763
rect -33 713 33 729
rect -15 691 15 713
rect -15 487 15 509
rect -33 471 33 487
rect -33 437 -17 471
rect 17 437 33 471
rect -33 421 33 437
rect -33 363 33 379
rect -33 329 -17 363
rect 17 329 33 363
rect -33 313 33 329
rect -15 291 15 313
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -313 15 -291
rect -33 -329 33 -313
rect -33 -363 -17 -329
rect 17 -363 33 -329
rect -33 -379 33 -363
rect -33 -437 33 -421
rect -33 -471 -17 -437
rect 17 -471 33 -437
rect -33 -487 33 -471
rect -15 -509 15 -487
rect -15 -713 15 -691
rect -33 -729 33 -713
rect -33 -763 -17 -729
rect 17 -763 33 -729
rect -33 -779 33 -763
rect -33 -837 33 -821
rect -33 -871 -17 -837
rect 17 -871 33 -837
rect -33 -887 33 -871
rect -15 -909 15 -887
rect -15 -1113 15 -1091
rect -33 -1129 33 -1113
rect -33 -1163 -17 -1129
rect 17 -1163 33 -1129
rect -33 -1179 33 -1163
rect -33 -1237 33 -1221
rect -33 -1271 -17 -1237
rect 17 -1271 33 -1237
rect -33 -1287 33 -1271
rect -15 -1309 15 -1287
rect -15 -1513 15 -1491
rect -33 -1529 33 -1513
rect -33 -1563 -17 -1529
rect 17 -1563 33 -1529
rect -33 -1579 33 -1563
<< polycont >>
rect -17 1529 17 1563
rect -17 1237 17 1271
rect -17 1129 17 1163
rect -17 837 17 871
rect -17 729 17 763
rect -17 437 17 471
rect -17 329 17 363
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -363 17 -329
rect -17 -471 17 -437
rect -17 -763 17 -729
rect -17 -871 17 -837
rect -17 -1163 17 -1129
rect -17 -1271 17 -1237
rect -17 -1563 17 -1529
<< locali >>
rect -33 1529 -17 1563
rect 17 1529 33 1563
rect -61 1479 -27 1495
rect -61 1305 -27 1321
rect 27 1479 61 1495
rect 27 1305 61 1321
rect -33 1237 -17 1271
rect 17 1237 33 1271
rect -33 1129 -17 1163
rect 17 1129 33 1163
rect -61 1079 -27 1095
rect -61 905 -27 921
rect 27 1079 61 1095
rect 27 905 61 921
rect -33 837 -17 871
rect 17 837 33 871
rect -33 729 -17 763
rect 17 729 33 763
rect -61 679 -27 695
rect -61 505 -27 521
rect 27 679 61 695
rect 27 505 61 521
rect -33 437 -17 471
rect 17 437 33 471
rect -33 329 -17 363
rect 17 329 33 363
rect -61 279 -27 295
rect -61 105 -27 121
rect 27 279 61 295
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -295 -27 -279
rect 27 -121 61 -105
rect 27 -295 61 -279
rect -33 -363 -17 -329
rect 17 -363 33 -329
rect -33 -471 -17 -437
rect 17 -471 33 -437
rect -61 -521 -27 -505
rect -61 -695 -27 -679
rect 27 -521 61 -505
rect 27 -695 61 -679
rect -33 -763 -17 -729
rect 17 -763 33 -729
rect -33 -871 -17 -837
rect 17 -871 33 -837
rect -61 -921 -27 -905
rect -61 -1095 -27 -1079
rect 27 -921 61 -905
rect 27 -1095 61 -1079
rect -33 -1163 -17 -1129
rect 17 -1163 33 -1129
rect -33 -1271 -17 -1237
rect 17 -1271 33 -1237
rect -61 -1321 -27 -1305
rect -61 -1495 -27 -1479
rect 27 -1321 61 -1305
rect 27 -1495 61 -1479
rect -33 -1563 -17 -1529
rect 17 -1563 33 -1529
<< viali >>
rect -17 1529 17 1563
rect -61 1321 -27 1479
rect 27 1321 61 1479
rect -17 1237 17 1271
rect -17 1129 17 1163
rect -61 921 -27 1079
rect 27 921 61 1079
rect -17 837 17 871
rect -17 729 17 763
rect -61 521 -27 679
rect 27 521 61 679
rect -17 437 17 471
rect -17 329 17 363
rect -61 121 -27 279
rect 27 121 61 279
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -279 -27 -121
rect 27 -279 61 -121
rect -17 -363 17 -329
rect -17 -471 17 -437
rect -61 -679 -27 -521
rect 27 -679 61 -521
rect -17 -763 17 -729
rect -17 -871 17 -837
rect -61 -1079 -27 -921
rect 27 -1079 61 -921
rect -17 -1163 17 -1129
rect -17 -1271 17 -1237
rect -61 -1479 -27 -1321
rect 27 -1479 61 -1321
rect -17 -1563 17 -1529
<< metal1 >>
rect -29 1563 29 1569
rect -29 1529 -17 1563
rect 17 1529 29 1563
rect -29 1523 29 1529
rect -67 1479 -21 1491
rect -67 1321 -61 1479
rect -27 1321 -21 1479
rect -67 1309 -21 1321
rect 21 1479 67 1491
rect 21 1321 27 1479
rect 61 1321 67 1479
rect 21 1309 67 1321
rect -29 1271 29 1277
rect -29 1237 -17 1271
rect 17 1237 29 1271
rect -29 1231 29 1237
rect -29 1163 29 1169
rect -29 1129 -17 1163
rect 17 1129 29 1163
rect -29 1123 29 1129
rect -67 1079 -21 1091
rect -67 921 -61 1079
rect -27 921 -21 1079
rect -67 909 -21 921
rect 21 1079 67 1091
rect 21 921 27 1079
rect 61 921 67 1079
rect 21 909 67 921
rect -29 871 29 877
rect -29 837 -17 871
rect 17 837 29 871
rect -29 831 29 837
rect -29 763 29 769
rect -29 729 -17 763
rect 17 729 29 763
rect -29 723 29 729
rect -67 679 -21 691
rect -67 521 -61 679
rect -27 521 -21 679
rect -67 509 -21 521
rect 21 679 67 691
rect 21 521 27 679
rect 61 521 67 679
rect 21 509 67 521
rect -29 471 29 477
rect -29 437 -17 471
rect 17 437 29 471
rect -29 431 29 437
rect -29 363 29 369
rect -29 329 -17 363
rect 17 329 29 363
rect -29 323 29 329
rect -67 279 -21 291
rect -67 121 -61 279
rect -27 121 -21 279
rect -67 109 -21 121
rect 21 279 67 291
rect 21 121 27 279
rect 61 121 67 279
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -279 -61 -121
rect -27 -279 -21 -121
rect -67 -291 -21 -279
rect 21 -121 67 -109
rect 21 -279 27 -121
rect 61 -279 67 -121
rect 21 -291 67 -279
rect -29 -329 29 -323
rect -29 -363 -17 -329
rect 17 -363 29 -329
rect -29 -369 29 -363
rect -29 -437 29 -431
rect -29 -471 -17 -437
rect 17 -471 29 -437
rect -29 -477 29 -471
rect -67 -521 -21 -509
rect -67 -679 -61 -521
rect -27 -679 -21 -521
rect -67 -691 -21 -679
rect 21 -521 67 -509
rect 21 -679 27 -521
rect 61 -679 67 -521
rect 21 -691 67 -679
rect -29 -729 29 -723
rect -29 -763 -17 -729
rect 17 -763 29 -729
rect -29 -769 29 -763
rect -29 -837 29 -831
rect -29 -871 -17 -837
rect 17 -871 29 -837
rect -29 -877 29 -871
rect -67 -921 -21 -909
rect -67 -1079 -61 -921
rect -27 -1079 -21 -921
rect -67 -1091 -21 -1079
rect 21 -921 67 -909
rect 21 -1079 27 -921
rect 61 -1079 67 -921
rect 21 -1091 67 -1079
rect -29 -1129 29 -1123
rect -29 -1163 -17 -1129
rect 17 -1163 29 -1129
rect -29 -1169 29 -1163
rect -29 -1237 29 -1231
rect -29 -1271 -17 -1237
rect 17 -1271 29 -1237
rect -29 -1277 29 -1271
rect -67 -1321 -21 -1309
rect -67 -1479 -61 -1321
rect -27 -1479 -21 -1321
rect -67 -1491 -21 -1479
rect 21 -1321 67 -1309
rect 21 -1479 27 -1321
rect 61 -1479 67 -1321
rect 21 -1491 67 -1479
rect -29 -1529 29 -1523
rect -29 -1563 -17 -1529
rect 17 -1563 29 -1529
rect -29 -1569 29 -1563
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 8 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
