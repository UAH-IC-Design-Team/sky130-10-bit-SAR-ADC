** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/tests/controller/controller_test.sch
**.subckt controller_test
V3 VDD GND 1.8V
V4 VSS GND 0
x1 VDD VSS sw_n_sp9 sw_n_sp8 sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2 sw_n_sp1 Gen_clk
+ reset_b sw_n8 sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 Vin_q sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6 sw_p_sp5
+ sw_p_sp4 sw_p_sp3 sw_p_sp2 sw_p_sp1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 bit10 bit9 bit8 bit7
+ bit6 bit5 bit4 bit3 bit2 bit1 done sw_sample controller
V1 clk GND PULSE 0 1.8V 10us 1ns 1ns 5us 10us
V5 reset_b GND PULSE 1.8V 0 5us 1ns 1ns 5us 1s
x2 VSS Vin_p VDD Vin_n Gen_clk clk Vin_q reset_b xor_clock_gen
V8 Vin_p GND PULSE 0 1.8V 10.1us 1ns 1ns 5us 20us
V9 Vin_n GND PULSE 0 1.8V 20.1us 1ns 1ns 5us 20us
**** begin user architecture code
 .lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


.options acct list
.temp 25
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
.control
tran 0.5u 200u
*plot RST_PLS clk+2 Pulse+4
plot done-4  sw_n_sp1 sw_n_sp2+2 sw_n_sp3+4 sw_n_sp4+6 sw_n_sp5+8 sw_n_sp6+10 sw_n_sp7+12
+ sw_n_sp8+14 sw_n_sp9+16 Vin_p+18 clk+20
plot done-4  sw_p_sp1 sw_p_sp2+2 sw_p_sp3+4 sw_p_sp4+6 sw_p_sp5+8 sw_p_sp6+10 sw_p_sp7+12
+ sw_p_sp8+14 sw_p_sp9+16 Vin_p+18 clk+20
plot done-4  sw_n1 sw_n2+2 sw_n3+4 sw_n4+6 sw_n5+8 sw_n6+10 sw_n7+12 sw_n8+14 Vin_p+16 clk+18
plot done-4  sw_p1 sw_p2+2 sw_p3+4 sw_p4+6 sw_p5+8 sw_p6+10 sw_p7+12 sw_p8+14 Vin_p+16 clk+18
plot done-4 bit1 bit2+2 bit3+4 bit4+6 bit5+8 bit6+10 bit7+12 bit8+14 bit9+16 bit10+18

plot done-4  sw_n_sp1 sw_n_sp2+2 sw_n_sp3+4 sw_n_sp4+6 sw_n_sp5+8 sw_n_sp6+10 sw_n_sp7+12
+ sw_n_sp8+14 sw_n_sp9+16 Vcmp+18 clk+20 sw_n1 sw_n2+2 sw_n3+4 sw_n4+6 sw_n5+8 sw_n6+10 sw_n7+12 sw_n8+14

plot done-4  sw_p_sp1 sw_p_sp2+2 sw_p_sp3+4 sw_p_sp4+6 sw_p_sp5+8 sw_p_sp6+10 sw_p_sp7+12
+ sw_p_sp8+14 sw_p_sp9+16 Vcmp+18 clk+20 sw_p1 sw_p2+2 sw_p3+4 sw_p4+6 sw_p5+8 sw_p6+10 sw_p7+12 sw_p8+14

plot clk reset_b+2 x1.cycle0+4 x1.cycle1+6 x1.cycle2+8 x1.cycle16+10 x1.cycle17+12 x1.cycle18+14
+ sw_sample+16 vin_p+18

plot reset_b-2 clk vin_p vin_n gen_clk
write controller_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  src/controller/controller.sym # of pins=12
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/controller/controller.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/controller/controller.sch
.subckt controller  VDD VSS sw_n_sp9 sw_n_sp8 sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2
+ sw_n_sp1 clk reset sw_n8 sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 Vcmp sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6
+ sw_p_sp5 sw_p_sp4 sw_p_sp3 sw_p_sp2 sw_p_sp1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 bit10 bit9 bit8
+ bit7 bit6 bit5 bit4 bit3 bit2 bit1 done sw_sample
*.ipin clk
*.opin sw_n_sp9,sw_n_sp8,sw_n_sp7,sw_n_sp6,sw_n_sp5,sw_n_sp4,sw_n_sp3,sw_n_sp2,sw_n_sp1
*.iopin VSS
*.iopin VDD
*.ipin reset
*.ipin Vcmp
*.opin sw_n8,sw_n7,sw_n6,sw_n5,sw_n4,sw_n3,sw_n2,sw_n1
*.opin sw_p_sp9,sw_p_sp8,sw_p_sp7,sw_p_sp6,sw_p_sp5,sw_p_sp4,sw_p_sp3,sw_p_sp2,sw_p_sp1
*.opin sw_p8,sw_p7,sw_p6,sw_p5,sw_p4,sw_p3,sw_p2,sw_p1
*.opin bit10,bit9,bit8,bit7,bit6,bit5,bit4,bit3,bit2,bit1
*.opin done
*.opin sw_sample
x95 cycle1 cycle2 cycle3 cycle4 VSS VSS VDD VDD net2 sky130_fd_sc_hd__or4_2
x96 cycle5 cycle6 cycle7 cycle8 VSS VSS VDD VDD net3 sky130_fd_sc_hd__or4_2
x97 cycle9 cycle10 cycle11 cycle12 VSS VSS VDD VDD net5 sky130_fd_sc_hd__or4_2
x2 clk clk_pulse VDD VSS reset pulse_generator
x3 VDD raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7 raw_bit6 raw_bit5 raw_bit4
+ raw_bit3 raw_bit2 raw_bit1 VSS reset bit10 bit9 bit8 bit7 bit6 bit5 bit4 bit3 bit2 bit1 done cycle31 dec
x4 raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7 raw_bit6 raw_bit5 raw_bit4
+ raw_bit3 raw_bit2 raw_bit1 cycle30 cycle29 cycle28 cycle27 cycle26 cycle25 cycle24 cycle23 cycle22 cycle21
+ cycle20 cycle19 cycle18 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 Vcmp net1 VDD VSS sw_n_sp9 sw_n_sp8
+ sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2 sw_n_sp1 sw_n8 sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2
+ sw_n1 sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6 sw_p_sp5 sw_p_sp4 sw_p_sp3 sw_p_sp2 sw_p_sp1 raw_bit_calculator
x1 clk VDD VSS clk_pulse reset cycle31 cycle30 cycle29 cycle28 cycle27 cycle26 cycle25 cycle24
+ cycle23 cycle22 cycle21 cycle20 cycle19 cycle18 cycle17 cycle16 cycle15 cycle14 cycle13 cycle12 cycle11
+ cycle10 cycle9 cycle8 cycle7 cycle6 cycle5 cycle4 cycle3 cycle2 cycle1 cycle0 shifted_clock_generator
x8 net2 net3 net5 net4 VSS VSS VDD VDD net6 sky130_fd_sc_hd__or4_2
x9 clk net6 reset VSS VSS VDD VDD sw_sample sky130_fd_sc_hd__dfrtn_1
x10 cycle13 cycle14 cycle15 VSS VSS VDD VDD net4 sky130_fd_sc_hd__or3_2
x6 cycle0 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x21 cycle2 net8 net7 VSS VSS VDD VDD Q_test1 sky130_fd_sc_hd__dfstp_1
x5 cycle0 VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_16
x7 Vcmp VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_16
XC1 VSS cycle2 sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=1 m=1
x11 cycle2 net10 net9 VSS VSS VDD VDD Q_test2 sky130_fd_sc_hd__dfstp_1
x12 cycle0 VSS VSS VDD VDD net9 sky130_fd_sc_hd__inv_16
x13 Vcmp VSS VSS VDD VDD net10 sky130_fd_sc_hd__inv_16
.ends


* expanding   symbol:  src/xor_clock_gen/xor_clock_gen.sym # of pins=8
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/xor_clock_gen/xor_clock_gen.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/xor_clock_gen/xor_clock_gen.sch
.subckt xor_clock_gen  VSS Vin_p VDD Vin_n Gen_clk Clk Vin_q Reset
*.ipin Vin_p
*.iopin VSS
*.opin Gen_clk
*.iopin VDD
*.ipin Vin_n
*.ipin Clk
*.ipin Reset
*.opin Vin_q
x1 Vin_p Vin_n VSS VSS VDD VDD net1 sky130_fd_sc_hd__xor2_1
x3 net1 VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
x6 net1 net2 Reset VSS VSS VDD VDD net5 net2 sky130_fd_sc_hd__dfrbp_1
x2 net7 net3 Reset VSS VSS VDD VDD net4 net3 sky130_fd_sc_hd__dfrbp_1
x4 net5 net4 VSS VSS VDD VDD net6 sky130_fd_sc_hd__xor2_1
x5 net6 VSS VSS VDD VDD net13 sky130_fd_sc_hd__inv_1
x7 net6 net8 Reset VSS VSS VDD VDD net11 net8 sky130_fd_sc_hd__dfrbp_1
x8 net13 net9 Reset VSS VSS VDD VDD net10 net9 sky130_fd_sc_hd__dfrbp_1
x9 net11 net10 VSS VSS VDD VDD net12 sky130_fd_sc_hd__xor2_1
x10 net12 VSS VSS VDD VDD net19 sky130_fd_sc_hd__inv_1
x11 net12 net14 Reset VSS VSS VDD VDD net17 net14 sky130_fd_sc_hd__dfrbp_1
x12 net19 net15 Reset VSS VSS VDD VDD net16 net15 sky130_fd_sc_hd__dfrbp_1
x13 net17 net16 VSS VSS VDD VDD net18 sky130_fd_sc_hd__xor2_1
x14 net6 Vin_p Reset VSS VSS VDD VDD net20 sky130_fd_sc_hd__dfrtp_1
x15 net18 VSS VSS VDD VDD net25 sky130_fd_sc_hd__inv_1
x16 net18 net21 Reset VSS VSS VDD VDD net24 net21 sky130_fd_sc_hd__dfrbp_1
x17 net25 net22 Reset VSS VSS VDD VDD net23 net22 sky130_fd_sc_hd__dfrbp_1
x18 net24 net23 VSS VSS VDD VDD Gen_clk sky130_fd_sc_hd__xor2_1
x19 net20 VSS VSS VDD VDD Vin_q sky130_fd_sc_hd__buf_16
.ends


* expanding   symbol:  src/pulse_generator/pulse_generator.sym # of pins=5
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/pulse_generator/pulse_generator.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/pulse_generator/pulse_generator.sch
.subckt pulse_generator  clk pulse VDD VSS RST_PLS
*.ipin clk
*.ipin RST_PLS
*.opin pulse
*.iopin VDD
*.iopin VSS
x1 clk net1 RST_PLS VSS VSS VDD VDD clk2 net1 sky130_fd_sc_hd__dfrbp_1
x2 clk2 net2 RST_PLS VSS VSS VDD VDD clk4 net2 sky130_fd_sc_hd__dfrbp_1
x3 clk4 net3 RST_PLS VSS VSS VDD VDD clk8 net3 sky130_fd_sc_hd__dfrbp_1
x4 clk8 net4 RST_PLS VSS VSS VDD VDD clk16 net4 sky130_fd_sc_hd__dfrbp_1
x5 delayed clk64 VSS VSS VDD VDD net7 sky130_fd_sc_hd__xor2_1
x9 clk16 net5 RST_PLS VSS VSS VDD VDD clk32 net5 sky130_fd_sc_hd__dfrbp_1
x10 clk32 net6 RST_PLS VSS VSS VDD VDD clk64 net6 sky130_fd_sc_hd__dfrbp_1
x6 clk clk64 RST_PLS VSS VSS VDD VDD delayed sky130_fd_sc_hd__dfrtp_1
x7 clk net7 RST_PLS VSS VSS VDD VDD pulse sky130_fd_sc_hd__dfrtn_1
.ends


* expanding   symbol:  src/dec/dec.sym # of pins=7
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/dec/dec.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/dec/dec.sch
.subckt dec  VDD raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7 raw_bit6
+ raw_bit5 raw_bit4 raw_bit3 raw_bit2 raw_bit1 VSS reset_b bit10 bit9 bit8 bit7 bit6 bit5 bit4 bit3 bit2 bit1
+ done dump_bus
*.iopin VDD
*.opin bit10,bit9,bit8,bit7,bit6,bit5,bit4,bit3,bit2,bit1
*.iopin VSS
*.ipin reset_b
*.ipin dump_bus
*.opin done
*.ipin
*+ raw_bit13,raw_bit12,raw_bit11,raw_bit10,raw_bit9,raw_bit8,raw_bit7,raw_bit6,raw_bit5,raw_bit4,raw_bit3,raw_bit2,raw_bit1
x62 raw_bit2 raw_bit1 net1 VSS VSS VDD VDD net16 net2 sky130_fd_sc_hd__fa_1
x64 raw_bit3 raw_bit1 net4 VSS VSS VDD VDD net1 net3 sky130_fd_sc_hd__fa_1
x67 dump_bus net2 reset_b VSS VSS VDD VDD bit2 sky130_fd_sc_hd__dfrtp_1
x68 dump_bus net3 reset_b VSS VSS VDD VDD bit3 sky130_fd_sc_hd__dfrtp_1
x65 raw_bit5 raw_bit4 net5 VSS VSS VDD VDD net4 net6 sky130_fd_sc_hd__fa_1
x69 raw_bit6 raw_bit4 net8 VSS VSS VDD VDD net5 net7 sky130_fd_sc_hd__fa_1
x70 dump_bus net6 reset_b VSS VSS VDD VDD bit4 sky130_fd_sc_hd__dfrtp_1
x71 dump_bus net7 reset_b VSS VSS VDD VDD bit5 sky130_fd_sc_hd__dfrtp_1
x72 raw_bit7 raw_bit4 net9 VSS VSS VDD VDD net8 net10 sky130_fd_sc_hd__fa_1
x73 raw_bit9 raw_bit8 net12 VSS VSS VDD VDD net9 net11 sky130_fd_sc_hd__fa_1
x74 dump_bus net10 reset_b VSS VSS VDD VDD bit6 sky130_fd_sc_hd__dfrtp_1
x75 dump_bus net11 reset_b VSS VSS VDD VDD bit7 sky130_fd_sc_hd__dfrtp_1
x76 raw_bit10 raw_bit8 net13 VSS VSS VDD VDD net12 net14 sky130_fd_sc_hd__fa_1
x77 raw_bit11 raw_bit8 raw_bit12 VSS VSS VDD VDD net13 net15 sky130_fd_sc_hd__fa_1
x78 dump_bus net14 reset_b VSS VSS VDD VDD bit8 sky130_fd_sc_hd__dfrtp_1
x79 dump_bus net15 reset_b VSS VSS VDD VDD bit9 sky130_fd_sc_hd__dfrtp_1
x80 dump_bus net16 reset_b VSS VSS VDD VDD bit1 sky130_fd_sc_hd__dfrtp_1
x81 dump_bus raw_bit13 reset_b VSS VSS VDD VDD bit10 sky130_fd_sc_hd__dfrtp_1
x82 dump_bus VSS VSS VDD VDD done sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  src/raw_bit_calculator/raw_bit_calculator.sym # of pins=10
** sym_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/raw_bit_calculator/raw_bit_calculator.sym
** sch_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/raw_bit_calculator/raw_bit_calculator.sch
.subckt raw_bit_calculator  raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7
+ raw_bit6 raw_bit5 raw_bit4 raw_bit3 raw_bit2 raw_bit1 cycle13 cycle12 cycle11 cycle10 cycle9 cycle8 cycle7
+ cycle6 cycle5 cycle4 cycle3 cycle2 cycle1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 Vcmp RESET VDD
+ VSS sw_n_sp9 sw_n_sp8 sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2 sw_n_sp1 sw_n8 sw_n7 sw_n6
+ sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6 sw_p_sp5 sw_p_sp4 sw_p_sp3 sw_p_sp2
+ sw_p_sp1
*.ipin
*+ cycle13,cycle12,cycle11,cycle10,cycle9,cycle8,cycle7,cycle6,cycle5,cycle4,cycle3,cycle2,cycle1
*.opin sw_n_sp9,sw_n_sp8,sw_n_sp7,sw_n_sp6,sw_n_sp5,sw_n_sp4,sw_n_sp3,sw_n_sp2,sw_n_sp1
*.iopin VSS
*.iopin VDD
*.opin sw_n8,sw_n7,sw_n6,sw_n5,sw_n4,sw_n3,sw_n2,sw_n1
*.opin sw_p_sp9,sw_p_sp8,sw_p_sp7,sw_p_sp6,sw_p_sp5,sw_p_sp4,sw_p_sp3,sw_p_sp2,sw_p_sp1
*.opin sw_p8,sw_p7,sw_p6,sw_p5,sw_p4,sw_p3,sw_p2,sw_p1
*.ipin Vcmp
*.ipin RESET
*.opin
*+ raw_bit13,raw_bit12,raw_bit11,raw_bit10,raw_bit9,raw_bit8,raw_bit7,raw_bit6,raw_bit5,raw_bit4,raw_bit3,raw_bit2,raw_bit1
x29 raw_bit1 Vcmp VSS VSS VDD VDD net50 sky130_fd_sc_hd__xor2_1
x31 raw_bit1 Vcmp VSS VSS VDD VDD net51 sky130_fd_sc_hd__xor2_1
x37 raw_bit4 Vcmp VSS VSS VDD VDD net52 sky130_fd_sc_hd__xor2_1
x40 raw_bit4 Vcmp VSS VSS VDD VDD net53 sky130_fd_sc_hd__xor2_1
x45 raw_bit4 Vcmp VSS VSS VDD VDD net54 sky130_fd_sc_hd__xor2_1
x100 cycle1 net10 net22 VSS VSS VDD VDD sw_p_sp1 sky130_fd_sc_hd__dfrtp_1
x99 Vcmp VSS VSS VDD VDD net10 sky130_fd_sc_hd__inv_1
x102 cycle1 Vcmp net22 VSS VSS VDD VDD sw_n_sp1 sky130_fd_sc_hd__dfrtp_1
x25 cycle1 Vcmp net24 VSS VSS VDD VDD sw_n_sp2 sky130_fd_sc_hd__dfrtp_1
x103 Vcmp VSS VSS VDD VDD net11 sky130_fd_sc_hd__inv_1
x104 cycle1 net11 net24 VSS VSS VDD VDD sw_p_sp2 sky130_fd_sc_hd__dfrtp_1
x21 net1 Vcmp RESET VSS VSS VDD VDD sw_n1 sky130_fd_sc_hd__dfstp_1
x22 net1 net12 RESET VSS VSS VDD VDD sw_p1 sky130_fd_sc_hd__dfstp_1
x105 Vcmp VSS VSS VDD VDD net12 sky130_fd_sc_hd__inv_1
x28 net3 Vcmp RESET VSS VSS VDD VDD sw_n2 sky130_fd_sc_hd__dfstp_1
x106 net3 net13 RESET VSS VSS VDD VDD sw_p2 sky130_fd_sc_hd__dfstp_1
x107 Vcmp VSS VSS VDD VDD net13 sky130_fd_sc_hd__inv_1
x109 Vcmp VSS VSS VDD VDD net14 sky130_fd_sc_hd__inv_1
x111 Vcmp VSS VSS VDD VDD net15 sky130_fd_sc_hd__inv_1
x27 cycle4 Vcmp net26 VSS VSS VDD VDD sw_n_sp3 sky130_fd_sc_hd__dfrtp_1
x35 cycle4 net14 net26 VSS VSS VDD VDD sw_p_sp3 sky130_fd_sc_hd__dfrtp_1
x41 cycle4 Vcmp net27 VSS VSS VDD VDD sw_n_sp4 sky130_fd_sc_hd__dfrtp_1
x108 cycle4 net15 net27 VSS VSS VDD VDD sw_p_sp4 sky130_fd_sc_hd__dfrtp_1
x110 cycle4 Vcmp net28 VSS VSS VDD VDD sw_n_sp5 sky130_fd_sc_hd__dfrtp_1
x112 cycle4 net16 net28 VSS VSS VDD VDD sw_p_sp5 sky130_fd_sc_hd__dfrtp_1
x113 Vcmp VSS VSS VDD VDD net16 sky130_fd_sc_hd__inv_1
x114 net5 net17 RESET VSS VSS VDD VDD sw_p3 sky130_fd_sc_hd__dfstp_1
x32 net5 Vcmp RESET VSS VSS VDD VDD sw_n3 sky130_fd_sc_hd__dfstp_1
x115 Vcmp VSS VSS VDD VDD net17 sky130_fd_sc_hd__inv_1
x38 net6 Vcmp RESET VSS VSS VDD VDD sw_n4 sky130_fd_sc_hd__dfstp_1
x116 net6 net18 RESET VSS VSS VDD VDD sw_p4 sky130_fd_sc_hd__dfstp_1
x117 Vcmp VSS VSS VDD VDD net18 sky130_fd_sc_hd__inv_1
x43 net7 Vcmp RESET VSS VSS VDD VDD sw_n5 sky130_fd_sc_hd__dfstp_1
x118 net7 net19 RESET VSS VSS VDD VDD sw_p5 sky130_fd_sc_hd__dfstp_1
x119 Vcmp VSS VSS VDD VDD net19 sky130_fd_sc_hd__inv_1
x132 cycle12 net20 RESET VSS VSS VDD VDD sw_p_sp9 sky130_fd_sc_hd__dfrtp_1
x133 Vcmp VSS VSS VDD VDD net20 sky130_fd_sc_hd__inv_1
x61 cycle12 Vcmp RESET VSS VSS VDD VDD sw_n_sp9 sky130_fd_sc_hd__dfrtp_1
x24 net50 VDD VSS net1 cycle2 net2 demux2
x30 net51 VDD VSS net3 cycle3 net4 demux2
x34 net52 VDD VSS net5 cycle5 net21 demux2
x39 net53 VDD VSS net6 cycle6 net8 demux2
x44 net54 VDD VSS net7 cycle7 net9 demux2
x1 net2 VSS VSS VDD VDD net23 sky130_fd_sc_hd__inv_1
x2 net4 VSS VSS VDD VDD net25 sky130_fd_sc_hd__inv_1
x3 cycle1 Vcmp RESET VSS VSS VDD VDD raw_bit1 sky130_fd_sc_hd__dfrtp_4
x4 cycle2 Vcmp RESET VSS VSS VDD VDD raw_bit2 sky130_fd_sc_hd__dfrtp_4
x5 cycle3 Vcmp RESET VSS VSS VDD VDD raw_bit3 sky130_fd_sc_hd__dfrtp_4
x6 cycle4 Vcmp RESET VSS VSS VDD VDD raw_bit4 sky130_fd_sc_hd__dfrtp_4
x7 cycle5 Vcmp RESET VSS VSS VDD VDD raw_bit5 sky130_fd_sc_hd__dfrtp_4
x8 cycle6 Vcmp RESET VSS VSS VDD VDD raw_bit6 sky130_fd_sc_hd__dfrtp_4
x9 cycle7 Vcmp RESET VSS VSS VDD VDD raw_bit7 sky130_fd_sc_hd__dfrtp_4
x10 cycle8 Vcmp RESET VSS VSS VDD VDD raw_bit8 sky130_fd_sc_hd__dfrtp_4
x11 cycle9 Vcmp RESET VSS VSS VDD VDD raw_bit9 sky130_fd_sc_hd__dfrtp_4
x12 cycle10 Vcmp RESET VSS VSS VDD VDD raw_bit10 sky130_fd_sc_hd__dfrtp_4
x13 cycle11 Vcmp RESET VSS VSS VDD VDD raw_bit11 sky130_fd_sc_hd__dfrtp_4
x14 cycle12 Vcmp RESET VSS VSS VDD VDD raw_bit12 sky130_fd_sc_hd__dfrtp_4
x15 cycle13 Vcmp RESET VSS VSS VDD VDD raw_bit13 sky130_fd_sc_hd__dfrtp_4
x18 net21 VSS VSS VDD VDD net29 sky130_fd_sc_hd__inv_1
x19 net8 VSS VSS VDD VDD net30 sky130_fd_sc_hd__inv_1
x20 net9 VSS VSS VDD VDD net31 sky130_fd_sc_hd__inv_1
x42 raw_bit8 Vcmp VSS VSS VDD VDD net55 sky130_fd_sc_hd__xor2_1
x62 raw_bit8 Vcmp VSS VSS VDD VDD net56 sky130_fd_sc_hd__xor2_1
x64 raw_bit8 Vcmp VSS VSS VDD VDD net57 sky130_fd_sc_hd__xor2_1
x65 Vcmp VSS VSS VDD VDD net37 sky130_fd_sc_hd__inv_1
x66 Vcmp VSS VSS VDD VDD net38 sky130_fd_sc_hd__inv_1
x67 cycle8 Vcmp net44 VSS VSS VDD VDD sw_n_sp6 sky130_fd_sc_hd__dfrtp_1
x68 cycle8 net37 net44 VSS VSS VDD VDD sw_p_sp6 sky130_fd_sc_hd__dfrtp_1
x69 cycle8 Vcmp net45 VSS VSS VDD VDD sw_n_sp7 sky130_fd_sc_hd__dfrtp_1
x70 cycle8 net38 net45 VSS VSS VDD VDD sw_p_sp7 sky130_fd_sc_hd__dfrtp_1
x71 cycle8 Vcmp net46 VSS VSS VDD VDD sw_n_sp8 sky130_fd_sc_hd__dfrtp_1
x72 cycle8 net39 net46 VSS VSS VDD VDD sw_p_sp8 sky130_fd_sc_hd__dfrtp_1
x73 Vcmp VSS VSS VDD VDD net39 sky130_fd_sc_hd__inv_1
x74 net32 net40 RESET VSS VSS VDD VDD sw_p6 sky130_fd_sc_hd__dfstp_1
x75 net32 Vcmp RESET VSS VSS VDD VDD sw_n6 sky130_fd_sc_hd__dfstp_1
x76 Vcmp VSS VSS VDD VDD net40 sky130_fd_sc_hd__inv_1
x77 net33 Vcmp RESET VSS VSS VDD VDD sw_n7 sky130_fd_sc_hd__dfstp_1
x78 net33 net41 RESET VSS VSS VDD VDD sw_p7 sky130_fd_sc_hd__dfstp_1
x79 Vcmp VSS VSS VDD VDD net41 sky130_fd_sc_hd__inv_1
x80 net34 Vcmp RESET VSS VSS VDD VDD sw_n8 sky130_fd_sc_hd__dfstp_1
x81 net34 net42 RESET VSS VSS VDD VDD sw_p8 sky130_fd_sc_hd__dfstp_1
x82 Vcmp VSS VSS VDD VDD net42 sky130_fd_sc_hd__inv_1
x83 net55 VDD VSS net32 cycle9 net43 demux2
x84 net56 VDD VSS net33 cycle10 net35 demux2
x85 net57 VDD VSS net34 cycle11 net36 demux2
x88 net43 VSS VSS VDD VDD net47 sky130_fd_sc_hd__inv_1
x89 net35 VSS VSS VDD VDD net48 sky130_fd_sc_hd__inv_1
x90 net36 VSS VSS VDD VDD net49 sky130_fd_sc_hd__inv_1
x46 net23 RESET VSS VSS VDD VDD net22 sky130_fd_sc_hd__and2_0
x23 net25 RESET VSS VSS VDD VDD net24 sky130_fd_sc_hd__and2_0
x26 net29 RESET VSS VSS VDD VDD net26 sky130_fd_sc_hd__and2_0
x16 net30 RESET VSS VSS VDD VDD net27 sky130_fd_sc_hd__and2_0
x17 net31 RESET VSS VSS VDD VDD net28 sky130_fd_sc_hd__and2_0
x33 net47 RESET VSS VSS VDD VDD net44 sky130_fd_sc_hd__and2_0
x36 net48 RESET VSS VSS VDD VDD net45 sky130_fd_sc_hd__and2_0
x47 net49 RESET VSS VSS VDD VDD net46 sky130_fd_sc_hd__and2_0
.ends


* expanding   symbol:  src/shifted_clock_generator/shifted_clock_generator.sym # of pins=6
** sym_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/shifted_clock_generator/shifted_clock_generator.sym
** sch_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/shifted_clock_generator/shifted_clock_generator.sch
.subckt shifted_clock_generator  clk VDD VSS clk_pulse reset_b cycle31 cycle30 cycle29 cycle28
+ cycle27 cycle26 cycle25 cycle24 cycle23 cycle22 cycle21 cycle20 cycle19 cycle18 cycle17 cycle16 cycle15
+ cycle14 cycle13 cycle12 cycle11 cycle10 cycle9 cycle8 cycle7 cycle6 cycle5 cycle4 cycle3 cycle2 cycle1
+ cycle0
*.ipin clk_pulse
*.opin
*+ cycle31,cycle30,cycle29,cycle28,cycle27,cycle26,cycle25,cycle24,cycle23,cycle22,cycle21,cycle20,cycle19,cycle18,cycle17,cycle16,cycle15,cycle14,cycle13,cycle12,cycle11,cycle10,cycle9,cycle8,cycle7,cycle6,cycle5,cycle4,cycle3,cycle2,cycle1,cycle0
*.iopin VSS
*.iopin VDD
*.ipin clk
*.ipin reset_b
x33 clk_pulse VSS VSS VDD VDD full_cycle0 sky130_fd_sc_hd__buf_12
x32 clk clk_pulse reset_b VSS VSS VDD VDD full_cycle1 sky130_fd_sc_hd__dfrtn_1
x1 clk full_cycle1 reset_b VSS VSS VDD VDD full_cycle2 sky130_fd_sc_hd__dfrtn_1
x2 clk full_cycle2 reset_b VSS VSS VDD VDD full_cycle3 sky130_fd_sc_hd__dfrtn_1
x3 clk full_cycle3 reset_b VSS VSS VDD VDD full_cycle4 sky130_fd_sc_hd__dfrtn_1
x4 clk full_cycle4 reset_b VSS VSS VDD VDD full_cycle5 sky130_fd_sc_hd__dfrtn_1
x5 clk full_cycle5 reset_b VSS VSS VDD VDD full_cycle6 sky130_fd_sc_hd__dfrtn_1
x6 clk full_cycle6 reset_b VSS VSS VDD VDD full_cycle7 sky130_fd_sc_hd__dfrtn_1
x7 clk full_cycle7 reset_b VSS VSS VDD VDD full_cycle8 sky130_fd_sc_hd__dfrtn_1
x8 clk full_cycle8 reset_b VSS VSS VDD VDD full_cycle9 sky130_fd_sc_hd__dfrtn_1
x9 clk full_cycle9 reset_b VSS VSS VDD VDD full_cycle10 sky130_fd_sc_hd__dfrtn_1
x10 clk full_cycle10 reset_b VSS VSS VDD VDD full_cycle11 sky130_fd_sc_hd__dfrtn_1
x11 clk full_cycle11 reset_b VSS VSS VDD VDD full_cycle12 sky130_fd_sc_hd__dfrtn_1
x12 clk full_cycle12 reset_b VSS VSS VDD VDD full_cycle13 sky130_fd_sc_hd__dfrtn_1
x13 clk full_cycle13 reset_b VSS VSS VDD VDD full_cycle14 sky130_fd_sc_hd__dfrtn_1
x14 clk full_cycle14 reset_b VSS VSS VDD VDD full_cycle15 sky130_fd_sc_hd__dfrtn_1
x15 clk full_cycle15 reset_b VSS VSS VDD VDD full_cycle16 sky130_fd_sc_hd__dfrtn_1
x16 clk full_cycle16 reset_b VSS VSS VDD VDD full_cycle17 sky130_fd_sc_hd__dfrtn_1
x17 clk full_cycle17 reset_b VSS VSS VDD VDD full_cycle18 sky130_fd_sc_hd__dfrtn_1
x18 clk full_cycle18 reset_b VSS VSS VDD VDD full_cycle19 sky130_fd_sc_hd__dfrtn_1
x19 clk full_cycle19 reset_b VSS VSS VDD VDD full_cycle20 sky130_fd_sc_hd__dfrtn_1
x20 clk full_cycle20 reset_b VSS VSS VDD VDD full_cycle21 sky130_fd_sc_hd__dfrtn_1
x21 clk full_cycle21 reset_b VSS VSS VDD VDD full_cycle22 sky130_fd_sc_hd__dfrtn_1
x22 clk full_cycle22 reset_b VSS VSS VDD VDD full_cycle23 sky130_fd_sc_hd__dfrtn_1
x23 clk full_cycle23 reset_b VSS VSS VDD VDD full_cycle24 sky130_fd_sc_hd__dfrtn_1
x24 clk full_cycle24 reset_b VSS VSS VDD VDD full_cycle25 sky130_fd_sc_hd__dfrtn_1
x25 clk full_cycle25 reset_b VSS VSS VDD VDD full_cycle26 sky130_fd_sc_hd__dfrtn_1
x26 clk full_cycle26 reset_b VSS VSS VDD VDD full_cycle27 sky130_fd_sc_hd__dfrtn_1
x27 clk full_cycle27 reset_b VSS VSS VDD VDD full_cycle28 sky130_fd_sc_hd__dfrtn_1
x28 clk full_cycle28 reset_b VSS VSS VDD VDD full_cycle29 sky130_fd_sc_hd__dfrtn_1
x29 clk full_cycle29 reset_b VSS VSS VDD VDD full_cycle30 sky130_fd_sc_hd__dfrtn_1
x30 clk full_cycle30 reset_b VSS VSS VDD VDD full_cycle31 sky130_fd_sc_hd__dfrtn_1
x35 clk full_cycle0 reset_b VSS VSS VDD VDD net1 sky130_fd_sc_hd__dfrtp_1
x36 net1 full_cycle0 VSS VSS VDD VDD net2 sky130_fd_sc_hd__and2_0
x39 clk full_cycle1 reset_b VSS VSS VDD VDD net3 sky130_fd_sc_hd__dfrtp_1
x40 net3 full_cycle1 VSS VSS VDD VDD net4 sky130_fd_sc_hd__and2_0
x31 clk full_cycle2 reset_b VSS VSS VDD VDD net5 sky130_fd_sc_hd__dfrtp_1
x34 net5 full_cycle2 VSS VSS VDD VDD net6 sky130_fd_sc_hd__and2_0
x37 clk full_cycle3 reset_b VSS VSS VDD VDD net7 sky130_fd_sc_hd__dfrtp_1
x38 net7 full_cycle3 VSS VSS VDD VDD cycle3 sky130_fd_sc_hd__and2_0
x41 clk full_cycle4 reset_b VSS VSS VDD VDD net8 sky130_fd_sc_hd__dfrtp_1
x42 net8 full_cycle4 VSS VSS VDD VDD cycle4 sky130_fd_sc_hd__and2_0
x43 clk full_cycle5 reset_b VSS VSS VDD VDD net9 sky130_fd_sc_hd__dfrtp_1
x44 net9 full_cycle5 VSS VSS VDD VDD cycle5 sky130_fd_sc_hd__and2_0
x45 clk full_cycle6 reset_b VSS VSS VDD VDD net10 sky130_fd_sc_hd__dfrtp_1
x46 net10 full_cycle6 VSS VSS VDD VDD cycle6 sky130_fd_sc_hd__and2_0
x47 clk full_cycle7 reset_b VSS VSS VDD VDD net11 sky130_fd_sc_hd__dfrtp_1
x48 net11 full_cycle7 VSS VSS VDD VDD cycle7 sky130_fd_sc_hd__and2_0
x49 clk full_cycle8 reset_b VSS VSS VDD VDD net12 sky130_fd_sc_hd__dfrtp_1
x50 net12 full_cycle8 VSS VSS VDD VDD cycle8 sky130_fd_sc_hd__and2_0
x51 clk full_cycle9 reset_b VSS VSS VDD VDD net13 sky130_fd_sc_hd__dfrtp_1
x52 net13 full_cycle9 VSS VSS VDD VDD cycle9 sky130_fd_sc_hd__and2_0
x53 clk full_cycle10 reset_b VSS VSS VDD VDD net14 sky130_fd_sc_hd__dfrtp_1
x54 net14 full_cycle10 VSS VSS VDD VDD cycle10 sky130_fd_sc_hd__and2_0
x55 clk full_cycle11 reset_b VSS VSS VDD VDD net15 sky130_fd_sc_hd__dfrtp_1
x56 net15 full_cycle11 VSS VSS VDD VDD cycle11 sky130_fd_sc_hd__and2_0
x57 clk full_cycle12 reset_b VSS VSS VDD VDD net16 sky130_fd_sc_hd__dfrtp_1
x58 net16 full_cycle12 VSS VSS VDD VDD cycle12 sky130_fd_sc_hd__and2_0
x59 clk full_cycle13 reset_b VSS VSS VDD VDD net17 sky130_fd_sc_hd__dfrtp_1
x60 net17 full_cycle13 VSS VSS VDD VDD cycle13 sky130_fd_sc_hd__and2_0
x61 clk full_cycle14 reset_b VSS VSS VDD VDD net18 sky130_fd_sc_hd__dfrtp_1
x62 net18 full_cycle14 VSS VSS VDD VDD cycle14 sky130_fd_sc_hd__and2_0
x63 clk full_cycle15 reset_b VSS VSS VDD VDD net19 sky130_fd_sc_hd__dfrtp_1
x64 net19 full_cycle15 VSS VSS VDD VDD cycle15 sky130_fd_sc_hd__and2_0
x65 clk full_cycle16 reset_b VSS VSS VDD VDD net20 sky130_fd_sc_hd__dfrtp_1
x66 net20 full_cycle16 VSS VSS VDD VDD cycle16 sky130_fd_sc_hd__and2_0
x67 clk full_cycle17 reset_b VSS VSS VDD VDD net21 sky130_fd_sc_hd__dfrtp_1
x68 net21 full_cycle17 VSS VSS VDD VDD cycle17 sky130_fd_sc_hd__and2_0
x69 clk full_cycle18 reset_b VSS VSS VDD VDD net22 sky130_fd_sc_hd__dfrtp_1
x70 net22 full_cycle18 VSS VSS VDD VDD cycle18 sky130_fd_sc_hd__and2_0
x71 clk full_cycle19 reset_b VSS VSS VDD VDD net23 sky130_fd_sc_hd__dfrtp_1
x72 net23 full_cycle19 VSS VSS VDD VDD cycle19 sky130_fd_sc_hd__and2_0
x73 clk full_cycle20 reset_b VSS VSS VDD VDD net24 sky130_fd_sc_hd__dfrtp_1
x74 net24 full_cycle20 VSS VSS VDD VDD cycle20 sky130_fd_sc_hd__and2_0
x75 clk full_cycle21 reset_b VSS VSS VDD VDD net25 sky130_fd_sc_hd__dfrtp_1
x76 net25 full_cycle21 VSS VSS VDD VDD cycle21 sky130_fd_sc_hd__and2_0
x77 clk full_cycle22 reset_b VSS VSS VDD VDD net26 sky130_fd_sc_hd__dfrtp_1
x78 net26 full_cycle22 VSS VSS VDD VDD cycle22 sky130_fd_sc_hd__and2_0
x79 clk full_cycle23 reset_b VSS VSS VDD VDD net27 sky130_fd_sc_hd__dfrtp_1
x80 net27 full_cycle23 VSS VSS VDD VDD cycle23 sky130_fd_sc_hd__and2_0
x81 clk full_cycle24 reset_b VSS VSS VDD VDD net28 sky130_fd_sc_hd__dfrtp_1
x82 net28 full_cycle24 VSS VSS VDD VDD cycle24 sky130_fd_sc_hd__and2_0
x83 clk full_cycle25 reset_b VSS VSS VDD VDD net29 sky130_fd_sc_hd__dfrtp_1
x84 net29 full_cycle25 VSS VSS VDD VDD cycle25 sky130_fd_sc_hd__and2_0
x85 clk full_cycle26 reset_b VSS VSS VDD VDD net30 sky130_fd_sc_hd__dfrtp_1
x86 net30 full_cycle26 VSS VSS VDD VDD cycle26 sky130_fd_sc_hd__and2_0
x87 clk full_cycle27 reset_b VSS VSS VDD VDD net31 sky130_fd_sc_hd__dfrtp_1
x88 net31 full_cycle27 VSS VSS VDD VDD cycle27 sky130_fd_sc_hd__and2_0
x89 clk full_cycle28 reset_b VSS VSS VDD VDD net32 sky130_fd_sc_hd__dfrtp_1
x90 net32 full_cycle28 VSS VSS VDD VDD cycle28 sky130_fd_sc_hd__and2_0
x91 clk full_cycle29 reset_b VSS VSS VDD VDD net33 sky130_fd_sc_hd__dfrtp_1
x92 net33 full_cycle29 VSS VSS VDD VDD cycle29 sky130_fd_sc_hd__and2_0
x93 clk full_cycle30 reset_b VSS VSS VDD VDD net34 sky130_fd_sc_hd__dfrtp_1
x94 net34 full_cycle30 VSS VSS VDD VDD cycle30 sky130_fd_sc_hd__and2_0
x95 clk full_cycle31 reset_b VSS VSS VDD VDD net35 sky130_fd_sc_hd__dfrtp_1
x96 net35 full_cycle31 VSS VSS VDD VDD cycle31 sky130_fd_sc_hd__and2_0
x97 net2 VSS VSS VDD VDD cycle0 sky130_fd_sc_hd__clkbuf_4
x98 net4 VSS VSS VDD VDD cycle1 sky130_fd_sc_hd__clkbuf_4
x99 net6 VSS VSS VDD VDD cycle2 sky130_fd_sc_hd__clkbuf_4
.ends


* expanding   symbol:  src/demux2/demux2.sym # of pins=6
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sch
.subckt demux2  S VDD VSS OUT_0 IN OUT_1
*.ipin S
*.opin OUT_0
*.ipin IN
*.opin OUT_1
*.iopin VDD
*.iopin VSS
x1 net1 IN VSS VSS VDD VDD OUT_0 sky130_fd_sc_hd__and2_0
x2 S IN VSS VSS VDD VDD OUT_1 sky130_fd_sc_hd__and2_0
x3 S VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_1
.ends

.GLOBAL GND
.end
