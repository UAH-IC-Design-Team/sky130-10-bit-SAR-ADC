magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< metal3 >>
rect -350 17962 349 17990
rect -350 13608 265 17962
rect 329 13608 349 17962
rect -350 13580 349 13608
rect -350 13452 349 13480
rect -350 9098 265 13452
rect 329 9098 349 13452
rect -350 9070 349 9098
rect -350 8942 349 8970
rect -350 4588 265 8942
rect 329 4588 349 8942
rect -350 4560 349 4588
rect -350 4432 349 4460
rect -350 78 265 4432
rect 329 78 349 4432
rect -350 50 349 78
rect -350 -78 349 -50
rect -350 -4432 265 -78
rect 329 -4432 349 -78
rect -350 -4460 349 -4432
rect -350 -4588 349 -4560
rect -350 -8942 265 -4588
rect 329 -8942 349 -4588
rect -350 -8970 349 -8942
rect -350 -9098 349 -9070
rect -350 -13452 265 -9098
rect 329 -13452 349 -9098
rect -350 -13480 349 -13452
rect -350 -13608 349 -13580
rect -350 -17962 265 -13608
rect 329 -17962 349 -13608
rect -350 -17990 349 -17962
<< via3 >>
rect 265 13608 329 17962
rect 265 9098 329 13452
rect 265 4588 329 8942
rect 265 78 329 4432
rect 265 -4432 329 -78
rect 265 -8942 329 -4588
rect 265 -13452 329 -9098
rect 265 -17962 329 -13608
<< mimcap >>
rect -250 17850 150 17890
rect -250 13720 -210 17850
rect 110 13720 150 17850
rect -250 13680 150 13720
rect -250 13340 150 13380
rect -250 9210 -210 13340
rect 110 9210 150 13340
rect -250 9170 150 9210
rect -250 8830 150 8870
rect -250 4700 -210 8830
rect 110 4700 150 8830
rect -250 4660 150 4700
rect -250 4320 150 4360
rect -250 190 -210 4320
rect 110 190 150 4320
rect -250 150 150 190
rect -250 -190 150 -150
rect -250 -4320 -210 -190
rect 110 -4320 150 -190
rect -250 -4360 150 -4320
rect -250 -4700 150 -4660
rect -250 -8830 -210 -4700
rect 110 -8830 150 -4700
rect -250 -8870 150 -8830
rect -250 -9210 150 -9170
rect -250 -13340 -210 -9210
rect 110 -13340 150 -9210
rect -250 -13380 150 -13340
rect -250 -13720 150 -13680
rect -250 -17850 -210 -13720
rect 110 -17850 150 -13720
rect -250 -17890 150 -17850
<< mimcapcontact >>
rect -210 13720 110 17850
rect -210 9210 110 13340
rect -210 4700 110 8830
rect -210 190 110 4320
rect -210 -4320 110 -190
rect -210 -8830 110 -4700
rect -210 -13340 110 -9210
rect -210 -17850 110 -13720
<< metal4 >>
rect -102 17851 2 18040
rect 218 17978 322 18040
rect 218 17962 345 17978
rect -211 17850 111 17851
rect -211 13720 -210 17850
rect 110 13720 111 17850
rect -211 13719 111 13720
rect -102 13341 2 13719
rect 218 13608 265 17962
rect 329 13608 345 17962
rect 218 13592 345 13608
rect 218 13468 322 13592
rect 218 13452 345 13468
rect -211 13340 111 13341
rect -211 9210 -210 13340
rect 110 9210 111 13340
rect -211 9209 111 9210
rect -102 8831 2 9209
rect 218 9098 265 13452
rect 329 9098 345 13452
rect 218 9082 345 9098
rect 218 8958 322 9082
rect 218 8942 345 8958
rect -211 8830 111 8831
rect -211 4700 -210 8830
rect 110 4700 111 8830
rect -211 4699 111 4700
rect -102 4321 2 4699
rect 218 4588 265 8942
rect 329 4588 345 8942
rect 218 4572 345 4588
rect 218 4448 322 4572
rect 218 4432 345 4448
rect -211 4320 111 4321
rect -211 190 -210 4320
rect 110 190 111 4320
rect -211 189 111 190
rect -102 -189 2 189
rect 218 78 265 4432
rect 329 78 345 4432
rect 218 62 345 78
rect 218 -62 322 62
rect 218 -78 345 -62
rect -211 -190 111 -189
rect -211 -4320 -210 -190
rect 110 -4320 111 -190
rect -211 -4321 111 -4320
rect -102 -4699 2 -4321
rect 218 -4432 265 -78
rect 329 -4432 345 -78
rect 218 -4448 345 -4432
rect 218 -4572 322 -4448
rect 218 -4588 345 -4572
rect -211 -4700 111 -4699
rect -211 -8830 -210 -4700
rect 110 -8830 111 -4700
rect -211 -8831 111 -8830
rect -102 -9209 2 -8831
rect 218 -8942 265 -4588
rect 329 -8942 345 -4588
rect 218 -8958 345 -8942
rect 218 -9082 322 -8958
rect 218 -9098 345 -9082
rect -211 -9210 111 -9209
rect -211 -13340 -210 -9210
rect 110 -13340 111 -9210
rect -211 -13341 111 -13340
rect -102 -13719 2 -13341
rect 218 -13452 265 -9098
rect 329 -13452 345 -9098
rect 218 -13468 345 -13452
rect 218 -13592 322 -13468
rect 218 -13608 345 -13592
rect -211 -13720 111 -13719
rect -211 -17850 -210 -13720
rect 110 -17850 111 -13720
rect -211 -17851 111 -17850
rect -102 -18040 2 -17851
rect 218 -17962 265 -13608
rect 329 -17962 345 -13608
rect 218 -17978 345 -17962
rect 218 -18040 322 -17978
<< properties >>
string FIXED_BBOX -350 13580 250 17990
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
