magic
tech sky130A
magscale 1 2
timestamp 1666819915
<< error_p >>
rect -29 -172 29 -166
rect -29 -206 -17 -172
rect -29 -212 29 -206
<< nwell >>
rect -109 -225 109 259
<< pmos >>
rect -15 -125 15 197
<< pdiff >>
rect -73 185 -15 197
rect -73 -113 -61 185
rect -27 -113 -15 185
rect -73 -125 -15 -113
rect 15 185 73 197
rect 15 -113 27 185
rect 61 -113 73 185
rect 15 -125 73 -113
<< pdiffc >>
rect -61 -113 -27 185
rect 27 -113 61 185
<< poly >>
rect -15 197 15 223
rect -15 -156 15 -125
rect -33 -172 33 -156
rect -33 -206 -17 -172
rect 17 -206 33 -172
rect -33 -222 33 -206
<< polycont >>
rect -17 -206 17 -172
<< locali >>
rect -61 185 -27 201
rect -61 -129 -27 -113
rect 27 185 61 201
rect 27 -129 61 -113
rect -33 -206 -17 -172
rect 17 -206 33 -172
<< viali >>
rect -61 -113 -27 185
rect 27 -16 61 88
rect -17 -206 17 -172
<< metal1 >>
rect -67 185 -21 197
rect -67 -113 -61 185
rect -27 -113 -21 185
rect 21 88 67 100
rect 21 -16 27 88
rect 61 -16 67 88
rect 21 -28 67 -16
rect -67 -125 -21 -113
rect -29 -172 29 -166
rect -29 -206 -17 -172
rect 17 -206 29 -172
rect -29 -212 29 -206
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 35 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
