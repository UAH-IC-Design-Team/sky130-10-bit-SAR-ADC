magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< error_p >>
rect -2227 139860 -2167 144270
rect -2147 139860 -2087 144270
rect -1508 139860 -1448 144270
rect -1428 139860 -1368 144270
rect -789 139860 -729 144270
rect -709 139860 -649 144270
rect -70 139860 -10 144270
rect 10 139860 70 144270
rect 649 139860 709 144270
rect 729 139860 789 144270
rect 1368 139860 1428 144270
rect 1448 139860 1508 144270
rect 2087 139860 2147 144270
rect 2167 139860 2227 144270
rect -2227 135350 -2167 139760
rect -2147 135350 -2087 139760
rect -1508 135350 -1448 139760
rect -1428 135350 -1368 139760
rect -789 135350 -729 139760
rect -709 135350 -649 139760
rect -70 135350 -10 139760
rect 10 135350 70 139760
rect 649 135350 709 139760
rect 729 135350 789 139760
rect 1368 135350 1428 139760
rect 1448 135350 1508 139760
rect 2087 135350 2147 139760
rect 2167 135350 2227 139760
rect -2227 130840 -2167 135250
rect -2147 130840 -2087 135250
rect -1508 130840 -1448 135250
rect -1428 130840 -1368 135250
rect -789 130840 -729 135250
rect -709 130840 -649 135250
rect -70 130840 -10 135250
rect 10 130840 70 135250
rect 649 130840 709 135250
rect 729 130840 789 135250
rect 1368 130840 1428 135250
rect 1448 130840 1508 135250
rect 2087 130840 2147 135250
rect 2167 130840 2227 135250
rect -2227 126330 -2167 130740
rect -2147 126330 -2087 130740
rect -1508 126330 -1448 130740
rect -1428 126330 -1368 130740
rect -789 126330 -729 130740
rect -709 126330 -649 130740
rect -70 126330 -10 130740
rect 10 126330 70 130740
rect 649 126330 709 130740
rect 729 126330 789 130740
rect 1368 126330 1428 130740
rect 1448 126330 1508 130740
rect 2087 126330 2147 130740
rect 2167 126330 2227 130740
rect -2227 121820 -2167 126230
rect -2147 121820 -2087 126230
rect -1508 121820 -1448 126230
rect -1428 121820 -1368 126230
rect -789 121820 -729 126230
rect -709 121820 -649 126230
rect -70 121820 -10 126230
rect 10 121820 70 126230
rect 649 121820 709 126230
rect 729 121820 789 126230
rect 1368 121820 1428 126230
rect 1448 121820 1508 126230
rect 2087 121820 2147 126230
rect 2167 121820 2227 126230
rect -2227 117310 -2167 121720
rect -2147 117310 -2087 121720
rect -1508 117310 -1448 121720
rect -1428 117310 -1368 121720
rect -789 117310 -729 121720
rect -709 117310 -649 121720
rect -70 117310 -10 121720
rect 10 117310 70 121720
rect 649 117310 709 121720
rect 729 117310 789 121720
rect 1368 117310 1428 121720
rect 1448 117310 1508 121720
rect 2087 117310 2147 121720
rect 2167 117310 2227 121720
rect -2227 112800 -2167 117210
rect -2147 112800 -2087 117210
rect -1508 112800 -1448 117210
rect -1428 112800 -1368 117210
rect -789 112800 -729 117210
rect -709 112800 -649 117210
rect -70 112800 -10 117210
rect 10 112800 70 117210
rect 649 112800 709 117210
rect 729 112800 789 117210
rect 1368 112800 1428 117210
rect 1448 112800 1508 117210
rect 2087 112800 2147 117210
rect 2167 112800 2227 117210
rect -2227 108290 -2167 112700
rect -2147 108290 -2087 112700
rect -1508 108290 -1448 112700
rect -1428 108290 -1368 112700
rect -789 108290 -729 112700
rect -709 108290 -649 112700
rect -70 108290 -10 112700
rect 10 108290 70 112700
rect 649 108290 709 112700
rect 729 108290 789 112700
rect 1368 108290 1428 112700
rect 1448 108290 1508 112700
rect 2087 108290 2147 112700
rect 2167 108290 2227 112700
rect -2227 103780 -2167 108190
rect -2147 103780 -2087 108190
rect -1508 103780 -1448 108190
rect -1428 103780 -1368 108190
rect -789 103780 -729 108190
rect -709 103780 -649 108190
rect -70 103780 -10 108190
rect 10 103780 70 108190
rect 649 103780 709 108190
rect 729 103780 789 108190
rect 1368 103780 1428 108190
rect 1448 103780 1508 108190
rect 2087 103780 2147 108190
rect 2167 103780 2227 108190
rect -2227 99270 -2167 103680
rect -2147 99270 -2087 103680
rect -1508 99270 -1448 103680
rect -1428 99270 -1368 103680
rect -789 99270 -729 103680
rect -709 99270 -649 103680
rect -70 99270 -10 103680
rect 10 99270 70 103680
rect 649 99270 709 103680
rect 729 99270 789 103680
rect 1368 99270 1428 103680
rect 1448 99270 1508 103680
rect 2087 99270 2147 103680
rect 2167 99270 2227 103680
rect -2227 94760 -2167 99170
rect -2147 94760 -2087 99170
rect -1508 94760 -1448 99170
rect -1428 94760 -1368 99170
rect -789 94760 -729 99170
rect -709 94760 -649 99170
rect -70 94760 -10 99170
rect 10 94760 70 99170
rect 649 94760 709 99170
rect 729 94760 789 99170
rect 1368 94760 1428 99170
rect 1448 94760 1508 99170
rect 2087 94760 2147 99170
rect 2167 94760 2227 99170
rect -2227 90250 -2167 94660
rect -2147 90250 -2087 94660
rect -1508 90250 -1448 94660
rect -1428 90250 -1368 94660
rect -789 90250 -729 94660
rect -709 90250 -649 94660
rect -70 90250 -10 94660
rect 10 90250 70 94660
rect 649 90250 709 94660
rect 729 90250 789 94660
rect 1368 90250 1428 94660
rect 1448 90250 1508 94660
rect 2087 90250 2147 94660
rect 2167 90250 2227 94660
rect -2227 85740 -2167 90150
rect -2147 85740 -2087 90150
rect -1508 85740 -1448 90150
rect -1428 85740 -1368 90150
rect -789 85740 -729 90150
rect -709 85740 -649 90150
rect -70 85740 -10 90150
rect 10 85740 70 90150
rect 649 85740 709 90150
rect 729 85740 789 90150
rect 1368 85740 1428 90150
rect 1448 85740 1508 90150
rect 2087 85740 2147 90150
rect 2167 85740 2227 90150
rect -2227 81230 -2167 85640
rect -2147 81230 -2087 85640
rect -1508 81230 -1448 85640
rect -1428 81230 -1368 85640
rect -789 81230 -729 85640
rect -709 81230 -649 85640
rect -70 81230 -10 85640
rect 10 81230 70 85640
rect 649 81230 709 85640
rect 729 81230 789 85640
rect 1368 81230 1428 85640
rect 1448 81230 1508 85640
rect 2087 81230 2147 85640
rect 2167 81230 2227 85640
rect -2227 76720 -2167 81130
rect -2147 76720 -2087 81130
rect -1508 76720 -1448 81130
rect -1428 76720 -1368 81130
rect -789 76720 -729 81130
rect -709 76720 -649 81130
rect -70 76720 -10 81130
rect 10 76720 70 81130
rect 649 76720 709 81130
rect 729 76720 789 81130
rect 1368 76720 1428 81130
rect 1448 76720 1508 81130
rect 2087 76720 2147 81130
rect 2167 76720 2227 81130
rect -2227 72210 -2167 76620
rect -2147 72210 -2087 76620
rect -1508 72210 -1448 76620
rect -1428 72210 -1368 76620
rect -789 72210 -729 76620
rect -709 72210 -649 76620
rect -70 72210 -10 76620
rect 10 72210 70 76620
rect 649 72210 709 76620
rect 729 72210 789 76620
rect 1368 72210 1428 76620
rect 1448 72210 1508 76620
rect 2087 72210 2147 76620
rect 2167 72210 2227 76620
rect -2227 67700 -2167 72110
rect -2147 67700 -2087 72110
rect -1508 67700 -1448 72110
rect -1428 67700 -1368 72110
rect -789 67700 -729 72110
rect -709 67700 -649 72110
rect -70 67700 -10 72110
rect 10 67700 70 72110
rect 649 67700 709 72110
rect 729 67700 789 72110
rect 1368 67700 1428 72110
rect 1448 67700 1508 72110
rect 2087 67700 2147 72110
rect 2167 67700 2227 72110
rect -2227 63190 -2167 67600
rect -2147 63190 -2087 67600
rect -1508 63190 -1448 67600
rect -1428 63190 -1368 67600
rect -789 63190 -729 67600
rect -709 63190 -649 67600
rect -70 63190 -10 67600
rect 10 63190 70 67600
rect 649 63190 709 67600
rect 729 63190 789 67600
rect 1368 63190 1428 67600
rect 1448 63190 1508 67600
rect 2087 63190 2147 67600
rect 2167 63190 2227 67600
rect -2227 58680 -2167 63090
rect -2147 58680 -2087 63090
rect -1508 58680 -1448 63090
rect -1428 58680 -1368 63090
rect -789 58680 -729 63090
rect -709 58680 -649 63090
rect -70 58680 -10 63090
rect 10 58680 70 63090
rect 649 58680 709 63090
rect 729 58680 789 63090
rect 1368 58680 1428 63090
rect 1448 58680 1508 63090
rect 2087 58680 2147 63090
rect 2167 58680 2227 63090
rect -2227 54170 -2167 58580
rect -2147 54170 -2087 58580
rect -1508 54170 -1448 58580
rect -1428 54170 -1368 58580
rect -789 54170 -729 58580
rect -709 54170 -649 58580
rect -70 54170 -10 58580
rect 10 54170 70 58580
rect 649 54170 709 58580
rect 729 54170 789 58580
rect 1368 54170 1428 58580
rect 1448 54170 1508 58580
rect 2087 54170 2147 58580
rect 2167 54170 2227 58580
rect -2227 49660 -2167 54070
rect -2147 49660 -2087 54070
rect -1508 49660 -1448 54070
rect -1428 49660 -1368 54070
rect -789 49660 -729 54070
rect -709 49660 -649 54070
rect -70 49660 -10 54070
rect 10 49660 70 54070
rect 649 49660 709 54070
rect 729 49660 789 54070
rect 1368 49660 1428 54070
rect 1448 49660 1508 54070
rect 2087 49660 2147 54070
rect 2167 49660 2227 54070
rect -2227 45150 -2167 49560
rect -2147 45150 -2087 49560
rect -1508 45150 -1448 49560
rect -1428 45150 -1368 49560
rect -789 45150 -729 49560
rect -709 45150 -649 49560
rect -70 45150 -10 49560
rect 10 45150 70 49560
rect 649 45150 709 49560
rect 729 45150 789 49560
rect 1368 45150 1428 49560
rect 1448 45150 1508 49560
rect 2087 45150 2147 49560
rect 2167 45150 2227 49560
rect -2227 40640 -2167 45050
rect -2147 40640 -2087 45050
rect -1508 40640 -1448 45050
rect -1428 40640 -1368 45050
rect -789 40640 -729 45050
rect -709 40640 -649 45050
rect -70 40640 -10 45050
rect 10 40640 70 45050
rect 649 40640 709 45050
rect 729 40640 789 45050
rect 1368 40640 1428 45050
rect 1448 40640 1508 45050
rect 2087 40640 2147 45050
rect 2167 40640 2227 45050
rect -2227 36130 -2167 40540
rect -2147 36130 -2087 40540
rect -1508 36130 -1448 40540
rect -1428 36130 -1368 40540
rect -789 36130 -729 40540
rect -709 36130 -649 40540
rect -70 36130 -10 40540
rect 10 36130 70 40540
rect 649 36130 709 40540
rect 729 36130 789 40540
rect 1368 36130 1428 40540
rect 1448 36130 1508 40540
rect 2087 36130 2147 40540
rect 2167 36130 2227 40540
rect -2227 31620 -2167 36030
rect -2147 31620 -2087 36030
rect -1508 31620 -1448 36030
rect -1428 31620 -1368 36030
rect -789 31620 -729 36030
rect -709 31620 -649 36030
rect -70 31620 -10 36030
rect 10 31620 70 36030
rect 649 31620 709 36030
rect 729 31620 789 36030
rect 1368 31620 1428 36030
rect 1448 31620 1508 36030
rect 2087 31620 2147 36030
rect 2167 31620 2227 36030
rect -2227 27110 -2167 31520
rect -2147 27110 -2087 31520
rect -1508 27110 -1448 31520
rect -1428 27110 -1368 31520
rect -789 27110 -729 31520
rect -709 27110 -649 31520
rect -70 27110 -10 31520
rect 10 27110 70 31520
rect 649 27110 709 31520
rect 729 27110 789 31520
rect 1368 27110 1428 31520
rect 1448 27110 1508 31520
rect 2087 27110 2147 31520
rect 2167 27110 2227 31520
rect -2227 22600 -2167 27010
rect -2147 22600 -2087 27010
rect -1508 22600 -1448 27010
rect -1428 22600 -1368 27010
rect -789 22600 -729 27010
rect -709 22600 -649 27010
rect -70 22600 -10 27010
rect 10 22600 70 27010
rect 649 22600 709 27010
rect 729 22600 789 27010
rect 1368 22600 1428 27010
rect 1448 22600 1508 27010
rect 2087 22600 2147 27010
rect 2167 22600 2227 27010
rect -2227 18090 -2167 22500
rect -2147 18090 -2087 22500
rect -1508 18090 -1448 22500
rect -1428 18090 -1368 22500
rect -789 18090 -729 22500
rect -709 18090 -649 22500
rect -70 18090 -10 22500
rect 10 18090 70 22500
rect 649 18090 709 22500
rect 729 18090 789 22500
rect 1368 18090 1428 22500
rect 1448 18090 1508 22500
rect 2087 18090 2147 22500
rect 2167 18090 2227 22500
rect -2227 13580 -2167 17990
rect -2147 13580 -2087 17990
rect -1508 13580 -1448 17990
rect -1428 13580 -1368 17990
rect -789 13580 -729 17990
rect -709 13580 -649 17990
rect -70 13580 -10 17990
rect 10 13580 70 17990
rect 649 13580 709 17990
rect 729 13580 789 17990
rect 1368 13580 1428 17990
rect 1448 13580 1508 17990
rect 2087 13580 2147 17990
rect 2167 13580 2227 17990
rect -2227 9070 -2167 13480
rect -2147 9070 -2087 13480
rect -1508 9070 -1448 13480
rect -1428 9070 -1368 13480
rect -789 9070 -729 13480
rect -709 9070 -649 13480
rect -70 9070 -10 13480
rect 10 9070 70 13480
rect 649 9070 709 13480
rect 729 9070 789 13480
rect 1368 9070 1428 13480
rect 1448 9070 1508 13480
rect 2087 9070 2147 13480
rect 2167 9070 2227 13480
rect -2227 4560 -2167 8970
rect -2147 4560 -2087 8970
rect -1508 4560 -1448 8970
rect -1428 4560 -1368 8970
rect -789 4560 -729 8970
rect -709 4560 -649 8970
rect -70 4560 -10 8970
rect 10 4560 70 8970
rect 649 4560 709 8970
rect 729 4560 789 8970
rect 1368 4560 1428 8970
rect 1448 4560 1508 8970
rect 2087 4560 2147 8970
rect 2167 4560 2227 8970
rect -2227 50 -2167 4460
rect -2147 50 -2087 4460
rect -1508 50 -1448 4460
rect -1428 50 -1368 4460
rect -789 50 -729 4460
rect -709 50 -649 4460
rect -70 50 -10 4460
rect 10 50 70 4460
rect 649 50 709 4460
rect 729 50 789 4460
rect 1368 50 1428 4460
rect 1448 50 1508 4460
rect 2087 50 2147 4460
rect 2167 50 2227 4460
rect -2227 -4460 -2167 -50
rect -2147 -4460 -2087 -50
rect -1508 -4460 -1448 -50
rect -1428 -4460 -1368 -50
rect -789 -4460 -729 -50
rect -709 -4460 -649 -50
rect -70 -4460 -10 -50
rect 10 -4460 70 -50
rect 649 -4460 709 -50
rect 729 -4460 789 -50
rect 1368 -4460 1428 -50
rect 1448 -4460 1508 -50
rect 2087 -4460 2147 -50
rect 2167 -4460 2227 -50
rect -2227 -8970 -2167 -4560
rect -2147 -8970 -2087 -4560
rect -1508 -8970 -1448 -4560
rect -1428 -8970 -1368 -4560
rect -789 -8970 -729 -4560
rect -709 -8970 -649 -4560
rect -70 -8970 -10 -4560
rect 10 -8970 70 -4560
rect 649 -8970 709 -4560
rect 729 -8970 789 -4560
rect 1368 -8970 1428 -4560
rect 1448 -8970 1508 -4560
rect 2087 -8970 2147 -4560
rect 2167 -8970 2227 -4560
rect -2227 -13480 -2167 -9070
rect -2147 -13480 -2087 -9070
rect -1508 -13480 -1448 -9070
rect -1428 -13480 -1368 -9070
rect -789 -13480 -729 -9070
rect -709 -13480 -649 -9070
rect -70 -13480 -10 -9070
rect 10 -13480 70 -9070
rect 649 -13480 709 -9070
rect 729 -13480 789 -9070
rect 1368 -13480 1428 -9070
rect 1448 -13480 1508 -9070
rect 2087 -13480 2147 -9070
rect 2167 -13480 2227 -9070
rect -2227 -17990 -2167 -13580
rect -2147 -17990 -2087 -13580
rect -1508 -17990 -1448 -13580
rect -1428 -17990 -1368 -13580
rect -789 -17990 -729 -13580
rect -709 -17990 -649 -13580
rect -70 -17990 -10 -13580
rect 10 -17990 70 -13580
rect 649 -17990 709 -13580
rect 729 -17990 789 -13580
rect 1368 -17990 1428 -13580
rect 1448 -17990 1508 -13580
rect 2087 -17990 2147 -13580
rect 2167 -17990 2227 -13580
rect -2227 -22500 -2167 -18090
rect -2147 -22500 -2087 -18090
rect -1508 -22500 -1448 -18090
rect -1428 -22500 -1368 -18090
rect -789 -22500 -729 -18090
rect -709 -22500 -649 -18090
rect -70 -22500 -10 -18090
rect 10 -22500 70 -18090
rect 649 -22500 709 -18090
rect 729 -22500 789 -18090
rect 1368 -22500 1428 -18090
rect 1448 -22500 1508 -18090
rect 2087 -22500 2147 -18090
rect 2167 -22500 2227 -18090
rect -2227 -27010 -2167 -22600
rect -2147 -27010 -2087 -22600
rect -1508 -27010 -1448 -22600
rect -1428 -27010 -1368 -22600
rect -789 -27010 -729 -22600
rect -709 -27010 -649 -22600
rect -70 -27010 -10 -22600
rect 10 -27010 70 -22600
rect 649 -27010 709 -22600
rect 729 -27010 789 -22600
rect 1368 -27010 1428 -22600
rect 1448 -27010 1508 -22600
rect 2087 -27010 2147 -22600
rect 2167 -27010 2227 -22600
rect -2227 -31520 -2167 -27110
rect -2147 -31520 -2087 -27110
rect -1508 -31520 -1448 -27110
rect -1428 -31520 -1368 -27110
rect -789 -31520 -729 -27110
rect -709 -31520 -649 -27110
rect -70 -31520 -10 -27110
rect 10 -31520 70 -27110
rect 649 -31520 709 -27110
rect 729 -31520 789 -27110
rect 1368 -31520 1428 -27110
rect 1448 -31520 1508 -27110
rect 2087 -31520 2147 -27110
rect 2167 -31520 2227 -27110
rect -2227 -36030 -2167 -31620
rect -2147 -36030 -2087 -31620
rect -1508 -36030 -1448 -31620
rect -1428 -36030 -1368 -31620
rect -789 -36030 -729 -31620
rect -709 -36030 -649 -31620
rect -70 -36030 -10 -31620
rect 10 -36030 70 -31620
rect 649 -36030 709 -31620
rect 729 -36030 789 -31620
rect 1368 -36030 1428 -31620
rect 1448 -36030 1508 -31620
rect 2087 -36030 2147 -31620
rect 2167 -36030 2227 -31620
rect -2227 -40540 -2167 -36130
rect -2147 -40540 -2087 -36130
rect -1508 -40540 -1448 -36130
rect -1428 -40540 -1368 -36130
rect -789 -40540 -729 -36130
rect -709 -40540 -649 -36130
rect -70 -40540 -10 -36130
rect 10 -40540 70 -36130
rect 649 -40540 709 -36130
rect 729 -40540 789 -36130
rect 1368 -40540 1428 -36130
rect 1448 -40540 1508 -36130
rect 2087 -40540 2147 -36130
rect 2167 -40540 2227 -36130
rect -2227 -45050 -2167 -40640
rect -2147 -45050 -2087 -40640
rect -1508 -45050 -1448 -40640
rect -1428 -45050 -1368 -40640
rect -789 -45050 -729 -40640
rect -709 -45050 -649 -40640
rect -70 -45050 -10 -40640
rect 10 -45050 70 -40640
rect 649 -45050 709 -40640
rect 729 -45050 789 -40640
rect 1368 -45050 1428 -40640
rect 1448 -45050 1508 -40640
rect 2087 -45050 2147 -40640
rect 2167 -45050 2227 -40640
rect -2227 -49560 -2167 -45150
rect -2147 -49560 -2087 -45150
rect -1508 -49560 -1448 -45150
rect -1428 -49560 -1368 -45150
rect -789 -49560 -729 -45150
rect -709 -49560 -649 -45150
rect -70 -49560 -10 -45150
rect 10 -49560 70 -45150
rect 649 -49560 709 -45150
rect 729 -49560 789 -45150
rect 1368 -49560 1428 -45150
rect 1448 -49560 1508 -45150
rect 2087 -49560 2147 -45150
rect 2167 -49560 2227 -45150
rect -2227 -54070 -2167 -49660
rect -2147 -54070 -2087 -49660
rect -1508 -54070 -1448 -49660
rect -1428 -54070 -1368 -49660
rect -789 -54070 -729 -49660
rect -709 -54070 -649 -49660
rect -70 -54070 -10 -49660
rect 10 -54070 70 -49660
rect 649 -54070 709 -49660
rect 729 -54070 789 -49660
rect 1368 -54070 1428 -49660
rect 1448 -54070 1508 -49660
rect 2087 -54070 2147 -49660
rect 2167 -54070 2227 -49660
rect -2227 -58580 -2167 -54170
rect -2147 -58580 -2087 -54170
rect -1508 -58580 -1448 -54170
rect -1428 -58580 -1368 -54170
rect -789 -58580 -729 -54170
rect -709 -58580 -649 -54170
rect -70 -58580 -10 -54170
rect 10 -58580 70 -54170
rect 649 -58580 709 -54170
rect 729 -58580 789 -54170
rect 1368 -58580 1428 -54170
rect 1448 -58580 1508 -54170
rect 2087 -58580 2147 -54170
rect 2167 -58580 2227 -54170
rect -2227 -63090 -2167 -58680
rect -2147 -63090 -2087 -58680
rect -1508 -63090 -1448 -58680
rect -1428 -63090 -1368 -58680
rect -789 -63090 -729 -58680
rect -709 -63090 -649 -58680
rect -70 -63090 -10 -58680
rect 10 -63090 70 -58680
rect 649 -63090 709 -58680
rect 729 -63090 789 -58680
rect 1368 -63090 1428 -58680
rect 1448 -63090 1508 -58680
rect 2087 -63090 2147 -58680
rect 2167 -63090 2227 -58680
rect -2227 -67600 -2167 -63190
rect -2147 -67600 -2087 -63190
rect -1508 -67600 -1448 -63190
rect -1428 -67600 -1368 -63190
rect -789 -67600 -729 -63190
rect -709 -67600 -649 -63190
rect -70 -67600 -10 -63190
rect 10 -67600 70 -63190
rect 649 -67600 709 -63190
rect 729 -67600 789 -63190
rect 1368 -67600 1428 -63190
rect 1448 -67600 1508 -63190
rect 2087 -67600 2147 -63190
rect 2167 -67600 2227 -63190
rect -2227 -72110 -2167 -67700
rect -2147 -72110 -2087 -67700
rect -1508 -72110 -1448 -67700
rect -1428 -72110 -1368 -67700
rect -789 -72110 -729 -67700
rect -709 -72110 -649 -67700
rect -70 -72110 -10 -67700
rect 10 -72110 70 -67700
rect 649 -72110 709 -67700
rect 729 -72110 789 -67700
rect 1368 -72110 1428 -67700
rect 1448 -72110 1508 -67700
rect 2087 -72110 2147 -67700
rect 2167 -72110 2227 -67700
rect -2227 -76620 -2167 -72210
rect -2147 -76620 -2087 -72210
rect -1508 -76620 -1448 -72210
rect -1428 -76620 -1368 -72210
rect -789 -76620 -729 -72210
rect -709 -76620 -649 -72210
rect -70 -76620 -10 -72210
rect 10 -76620 70 -72210
rect 649 -76620 709 -72210
rect 729 -76620 789 -72210
rect 1368 -76620 1428 -72210
rect 1448 -76620 1508 -72210
rect 2087 -76620 2147 -72210
rect 2167 -76620 2227 -72210
rect -2227 -81130 -2167 -76720
rect -2147 -81130 -2087 -76720
rect -1508 -81130 -1448 -76720
rect -1428 -81130 -1368 -76720
rect -789 -81130 -729 -76720
rect -709 -81130 -649 -76720
rect -70 -81130 -10 -76720
rect 10 -81130 70 -76720
rect 649 -81130 709 -76720
rect 729 -81130 789 -76720
rect 1368 -81130 1428 -76720
rect 1448 -81130 1508 -76720
rect 2087 -81130 2147 -76720
rect 2167 -81130 2227 -76720
rect -2227 -85640 -2167 -81230
rect -2147 -85640 -2087 -81230
rect -1508 -85640 -1448 -81230
rect -1428 -85640 -1368 -81230
rect -789 -85640 -729 -81230
rect -709 -85640 -649 -81230
rect -70 -85640 -10 -81230
rect 10 -85640 70 -81230
rect 649 -85640 709 -81230
rect 729 -85640 789 -81230
rect 1368 -85640 1428 -81230
rect 1448 -85640 1508 -81230
rect 2087 -85640 2147 -81230
rect 2167 -85640 2227 -81230
rect -2227 -90150 -2167 -85740
rect -2147 -90150 -2087 -85740
rect -1508 -90150 -1448 -85740
rect -1428 -90150 -1368 -85740
rect -789 -90150 -729 -85740
rect -709 -90150 -649 -85740
rect -70 -90150 -10 -85740
rect 10 -90150 70 -85740
rect 649 -90150 709 -85740
rect 729 -90150 789 -85740
rect 1368 -90150 1428 -85740
rect 1448 -90150 1508 -85740
rect 2087 -90150 2147 -85740
rect 2167 -90150 2227 -85740
rect -2227 -94660 -2167 -90250
rect -2147 -94660 -2087 -90250
rect -1508 -94660 -1448 -90250
rect -1428 -94660 -1368 -90250
rect -789 -94660 -729 -90250
rect -709 -94660 -649 -90250
rect -70 -94660 -10 -90250
rect 10 -94660 70 -90250
rect 649 -94660 709 -90250
rect 729 -94660 789 -90250
rect 1368 -94660 1428 -90250
rect 1448 -94660 1508 -90250
rect 2087 -94660 2147 -90250
rect 2167 -94660 2227 -90250
rect -2227 -99170 -2167 -94760
rect -2147 -99170 -2087 -94760
rect -1508 -99170 -1448 -94760
rect -1428 -99170 -1368 -94760
rect -789 -99170 -729 -94760
rect -709 -99170 -649 -94760
rect -70 -99170 -10 -94760
rect 10 -99170 70 -94760
rect 649 -99170 709 -94760
rect 729 -99170 789 -94760
rect 1368 -99170 1428 -94760
rect 1448 -99170 1508 -94760
rect 2087 -99170 2147 -94760
rect 2167 -99170 2227 -94760
rect -2227 -103680 -2167 -99270
rect -2147 -103680 -2087 -99270
rect -1508 -103680 -1448 -99270
rect -1428 -103680 -1368 -99270
rect -789 -103680 -729 -99270
rect -709 -103680 -649 -99270
rect -70 -103680 -10 -99270
rect 10 -103680 70 -99270
rect 649 -103680 709 -99270
rect 729 -103680 789 -99270
rect 1368 -103680 1428 -99270
rect 1448 -103680 1508 -99270
rect 2087 -103680 2147 -99270
rect 2167 -103680 2227 -99270
rect -2227 -108190 -2167 -103780
rect -2147 -108190 -2087 -103780
rect -1508 -108190 -1448 -103780
rect -1428 -108190 -1368 -103780
rect -789 -108190 -729 -103780
rect -709 -108190 -649 -103780
rect -70 -108190 -10 -103780
rect 10 -108190 70 -103780
rect 649 -108190 709 -103780
rect 729 -108190 789 -103780
rect 1368 -108190 1428 -103780
rect 1448 -108190 1508 -103780
rect 2087 -108190 2147 -103780
rect 2167 -108190 2227 -103780
rect -2227 -112700 -2167 -108290
rect -2147 -112700 -2087 -108290
rect -1508 -112700 -1448 -108290
rect -1428 -112700 -1368 -108290
rect -789 -112700 -729 -108290
rect -709 -112700 -649 -108290
rect -70 -112700 -10 -108290
rect 10 -112700 70 -108290
rect 649 -112700 709 -108290
rect 729 -112700 789 -108290
rect 1368 -112700 1428 -108290
rect 1448 -112700 1508 -108290
rect 2087 -112700 2147 -108290
rect 2167 -112700 2227 -108290
rect -2227 -117210 -2167 -112800
rect -2147 -117210 -2087 -112800
rect -1508 -117210 -1448 -112800
rect -1428 -117210 -1368 -112800
rect -789 -117210 -729 -112800
rect -709 -117210 -649 -112800
rect -70 -117210 -10 -112800
rect 10 -117210 70 -112800
rect 649 -117210 709 -112800
rect 729 -117210 789 -112800
rect 1368 -117210 1428 -112800
rect 1448 -117210 1508 -112800
rect 2087 -117210 2147 -112800
rect 2167 -117210 2227 -112800
rect -2227 -121720 -2167 -117310
rect -2147 -121720 -2087 -117310
rect -1508 -121720 -1448 -117310
rect -1428 -121720 -1368 -117310
rect -789 -121720 -729 -117310
rect -709 -121720 -649 -117310
rect -70 -121720 -10 -117310
rect 10 -121720 70 -117310
rect 649 -121720 709 -117310
rect 729 -121720 789 -117310
rect 1368 -121720 1428 -117310
rect 1448 -121720 1508 -117310
rect 2087 -121720 2147 -117310
rect 2167 -121720 2227 -117310
rect -2227 -126230 -2167 -121820
rect -2147 -126230 -2087 -121820
rect -1508 -126230 -1448 -121820
rect -1428 -126230 -1368 -121820
rect -789 -126230 -729 -121820
rect -709 -126230 -649 -121820
rect -70 -126230 -10 -121820
rect 10 -126230 70 -121820
rect 649 -126230 709 -121820
rect 729 -126230 789 -121820
rect 1368 -126230 1428 -121820
rect 1448 -126230 1508 -121820
rect 2087 -126230 2147 -121820
rect 2167 -126230 2227 -121820
rect -2227 -130740 -2167 -126330
rect -2147 -130740 -2087 -126330
rect -1508 -130740 -1448 -126330
rect -1428 -130740 -1368 -126330
rect -789 -130740 -729 -126330
rect -709 -130740 -649 -126330
rect -70 -130740 -10 -126330
rect 10 -130740 70 -126330
rect 649 -130740 709 -126330
rect 729 -130740 789 -126330
rect 1368 -130740 1428 -126330
rect 1448 -130740 1508 -126330
rect 2087 -130740 2147 -126330
rect 2167 -130740 2227 -126330
rect -2227 -135250 -2167 -130840
rect -2147 -135250 -2087 -130840
rect -1508 -135250 -1448 -130840
rect -1428 -135250 -1368 -130840
rect -789 -135250 -729 -130840
rect -709 -135250 -649 -130840
rect -70 -135250 -10 -130840
rect 10 -135250 70 -130840
rect 649 -135250 709 -130840
rect 729 -135250 789 -130840
rect 1368 -135250 1428 -130840
rect 1448 -135250 1508 -130840
rect 2087 -135250 2147 -130840
rect 2167 -135250 2227 -130840
rect -2227 -139760 -2167 -135350
rect -2147 -139760 -2087 -135350
rect -1508 -139760 -1448 -135350
rect -1428 -139760 -1368 -135350
rect -789 -139760 -729 -135350
rect -709 -139760 -649 -135350
rect -70 -139760 -10 -135350
rect 10 -139760 70 -135350
rect 649 -139760 709 -135350
rect 729 -139760 789 -135350
rect 1368 -139760 1428 -135350
rect 1448 -139760 1508 -135350
rect 2087 -139760 2147 -135350
rect 2167 -139760 2227 -135350
rect -2227 -144270 -2167 -139860
rect -2147 -144270 -2087 -139860
rect -1508 -144270 -1448 -139860
rect -1428 -144270 -1368 -139860
rect -789 -144270 -729 -139860
rect -709 -144270 -649 -139860
rect -70 -144270 -10 -139860
rect 10 -144270 70 -139860
rect 649 -144270 709 -139860
rect 729 -144270 789 -139860
rect 1368 -144270 1428 -139860
rect 1448 -144270 1508 -139860
rect 2087 -144270 2147 -139860
rect 2167 -144270 2227 -139860
<< metal3 >>
rect -2866 144242 -2167 144270
rect -2866 139888 -2251 144242
rect -2187 139888 -2167 144242
rect -2866 139860 -2167 139888
rect -2147 144242 -1448 144270
rect -2147 139888 -1532 144242
rect -1468 139888 -1448 144242
rect -2147 139860 -1448 139888
rect -1428 144242 -729 144270
rect -1428 139888 -813 144242
rect -749 139888 -729 144242
rect -1428 139860 -729 139888
rect -709 144242 -10 144270
rect -709 139888 -94 144242
rect -30 139888 -10 144242
rect -709 139860 -10 139888
rect 10 144242 709 144270
rect 10 139888 625 144242
rect 689 139888 709 144242
rect 10 139860 709 139888
rect 729 144242 1428 144270
rect 729 139888 1344 144242
rect 1408 139888 1428 144242
rect 729 139860 1428 139888
rect 1448 144242 2147 144270
rect 1448 139888 2063 144242
rect 2127 139888 2147 144242
rect 1448 139860 2147 139888
rect 2167 144242 2866 144270
rect 2167 139888 2782 144242
rect 2846 139888 2866 144242
rect 2167 139860 2866 139888
rect -2866 139732 -2167 139760
rect -2866 135378 -2251 139732
rect -2187 135378 -2167 139732
rect -2866 135350 -2167 135378
rect -2147 139732 -1448 139760
rect -2147 135378 -1532 139732
rect -1468 135378 -1448 139732
rect -2147 135350 -1448 135378
rect -1428 139732 -729 139760
rect -1428 135378 -813 139732
rect -749 135378 -729 139732
rect -1428 135350 -729 135378
rect -709 139732 -10 139760
rect -709 135378 -94 139732
rect -30 135378 -10 139732
rect -709 135350 -10 135378
rect 10 139732 709 139760
rect 10 135378 625 139732
rect 689 135378 709 139732
rect 10 135350 709 135378
rect 729 139732 1428 139760
rect 729 135378 1344 139732
rect 1408 135378 1428 139732
rect 729 135350 1428 135378
rect 1448 139732 2147 139760
rect 1448 135378 2063 139732
rect 2127 135378 2147 139732
rect 1448 135350 2147 135378
rect 2167 139732 2866 139760
rect 2167 135378 2782 139732
rect 2846 135378 2866 139732
rect 2167 135350 2866 135378
rect -2866 135222 -2167 135250
rect -2866 130868 -2251 135222
rect -2187 130868 -2167 135222
rect -2866 130840 -2167 130868
rect -2147 135222 -1448 135250
rect -2147 130868 -1532 135222
rect -1468 130868 -1448 135222
rect -2147 130840 -1448 130868
rect -1428 135222 -729 135250
rect -1428 130868 -813 135222
rect -749 130868 -729 135222
rect -1428 130840 -729 130868
rect -709 135222 -10 135250
rect -709 130868 -94 135222
rect -30 130868 -10 135222
rect -709 130840 -10 130868
rect 10 135222 709 135250
rect 10 130868 625 135222
rect 689 130868 709 135222
rect 10 130840 709 130868
rect 729 135222 1428 135250
rect 729 130868 1344 135222
rect 1408 130868 1428 135222
rect 729 130840 1428 130868
rect 1448 135222 2147 135250
rect 1448 130868 2063 135222
rect 2127 130868 2147 135222
rect 1448 130840 2147 130868
rect 2167 135222 2866 135250
rect 2167 130868 2782 135222
rect 2846 130868 2866 135222
rect 2167 130840 2866 130868
rect -2866 130712 -2167 130740
rect -2866 126358 -2251 130712
rect -2187 126358 -2167 130712
rect -2866 126330 -2167 126358
rect -2147 130712 -1448 130740
rect -2147 126358 -1532 130712
rect -1468 126358 -1448 130712
rect -2147 126330 -1448 126358
rect -1428 130712 -729 130740
rect -1428 126358 -813 130712
rect -749 126358 -729 130712
rect -1428 126330 -729 126358
rect -709 130712 -10 130740
rect -709 126358 -94 130712
rect -30 126358 -10 130712
rect -709 126330 -10 126358
rect 10 130712 709 130740
rect 10 126358 625 130712
rect 689 126358 709 130712
rect 10 126330 709 126358
rect 729 130712 1428 130740
rect 729 126358 1344 130712
rect 1408 126358 1428 130712
rect 729 126330 1428 126358
rect 1448 130712 2147 130740
rect 1448 126358 2063 130712
rect 2127 126358 2147 130712
rect 1448 126330 2147 126358
rect 2167 130712 2866 130740
rect 2167 126358 2782 130712
rect 2846 126358 2866 130712
rect 2167 126330 2866 126358
rect -2866 126202 -2167 126230
rect -2866 121848 -2251 126202
rect -2187 121848 -2167 126202
rect -2866 121820 -2167 121848
rect -2147 126202 -1448 126230
rect -2147 121848 -1532 126202
rect -1468 121848 -1448 126202
rect -2147 121820 -1448 121848
rect -1428 126202 -729 126230
rect -1428 121848 -813 126202
rect -749 121848 -729 126202
rect -1428 121820 -729 121848
rect -709 126202 -10 126230
rect -709 121848 -94 126202
rect -30 121848 -10 126202
rect -709 121820 -10 121848
rect 10 126202 709 126230
rect 10 121848 625 126202
rect 689 121848 709 126202
rect 10 121820 709 121848
rect 729 126202 1428 126230
rect 729 121848 1344 126202
rect 1408 121848 1428 126202
rect 729 121820 1428 121848
rect 1448 126202 2147 126230
rect 1448 121848 2063 126202
rect 2127 121848 2147 126202
rect 1448 121820 2147 121848
rect 2167 126202 2866 126230
rect 2167 121848 2782 126202
rect 2846 121848 2866 126202
rect 2167 121820 2866 121848
rect -2866 121692 -2167 121720
rect -2866 117338 -2251 121692
rect -2187 117338 -2167 121692
rect -2866 117310 -2167 117338
rect -2147 121692 -1448 121720
rect -2147 117338 -1532 121692
rect -1468 117338 -1448 121692
rect -2147 117310 -1448 117338
rect -1428 121692 -729 121720
rect -1428 117338 -813 121692
rect -749 117338 -729 121692
rect -1428 117310 -729 117338
rect -709 121692 -10 121720
rect -709 117338 -94 121692
rect -30 117338 -10 121692
rect -709 117310 -10 117338
rect 10 121692 709 121720
rect 10 117338 625 121692
rect 689 117338 709 121692
rect 10 117310 709 117338
rect 729 121692 1428 121720
rect 729 117338 1344 121692
rect 1408 117338 1428 121692
rect 729 117310 1428 117338
rect 1448 121692 2147 121720
rect 1448 117338 2063 121692
rect 2127 117338 2147 121692
rect 1448 117310 2147 117338
rect 2167 121692 2866 121720
rect 2167 117338 2782 121692
rect 2846 117338 2866 121692
rect 2167 117310 2866 117338
rect -2866 117182 -2167 117210
rect -2866 112828 -2251 117182
rect -2187 112828 -2167 117182
rect -2866 112800 -2167 112828
rect -2147 117182 -1448 117210
rect -2147 112828 -1532 117182
rect -1468 112828 -1448 117182
rect -2147 112800 -1448 112828
rect -1428 117182 -729 117210
rect -1428 112828 -813 117182
rect -749 112828 -729 117182
rect -1428 112800 -729 112828
rect -709 117182 -10 117210
rect -709 112828 -94 117182
rect -30 112828 -10 117182
rect -709 112800 -10 112828
rect 10 117182 709 117210
rect 10 112828 625 117182
rect 689 112828 709 117182
rect 10 112800 709 112828
rect 729 117182 1428 117210
rect 729 112828 1344 117182
rect 1408 112828 1428 117182
rect 729 112800 1428 112828
rect 1448 117182 2147 117210
rect 1448 112828 2063 117182
rect 2127 112828 2147 117182
rect 1448 112800 2147 112828
rect 2167 117182 2866 117210
rect 2167 112828 2782 117182
rect 2846 112828 2866 117182
rect 2167 112800 2866 112828
rect -2866 112672 -2167 112700
rect -2866 108318 -2251 112672
rect -2187 108318 -2167 112672
rect -2866 108290 -2167 108318
rect -2147 112672 -1448 112700
rect -2147 108318 -1532 112672
rect -1468 108318 -1448 112672
rect -2147 108290 -1448 108318
rect -1428 112672 -729 112700
rect -1428 108318 -813 112672
rect -749 108318 -729 112672
rect -1428 108290 -729 108318
rect -709 112672 -10 112700
rect -709 108318 -94 112672
rect -30 108318 -10 112672
rect -709 108290 -10 108318
rect 10 112672 709 112700
rect 10 108318 625 112672
rect 689 108318 709 112672
rect 10 108290 709 108318
rect 729 112672 1428 112700
rect 729 108318 1344 112672
rect 1408 108318 1428 112672
rect 729 108290 1428 108318
rect 1448 112672 2147 112700
rect 1448 108318 2063 112672
rect 2127 108318 2147 112672
rect 1448 108290 2147 108318
rect 2167 112672 2866 112700
rect 2167 108318 2782 112672
rect 2846 108318 2866 112672
rect 2167 108290 2866 108318
rect -2866 108162 -2167 108190
rect -2866 103808 -2251 108162
rect -2187 103808 -2167 108162
rect -2866 103780 -2167 103808
rect -2147 108162 -1448 108190
rect -2147 103808 -1532 108162
rect -1468 103808 -1448 108162
rect -2147 103780 -1448 103808
rect -1428 108162 -729 108190
rect -1428 103808 -813 108162
rect -749 103808 -729 108162
rect -1428 103780 -729 103808
rect -709 108162 -10 108190
rect -709 103808 -94 108162
rect -30 103808 -10 108162
rect -709 103780 -10 103808
rect 10 108162 709 108190
rect 10 103808 625 108162
rect 689 103808 709 108162
rect 10 103780 709 103808
rect 729 108162 1428 108190
rect 729 103808 1344 108162
rect 1408 103808 1428 108162
rect 729 103780 1428 103808
rect 1448 108162 2147 108190
rect 1448 103808 2063 108162
rect 2127 103808 2147 108162
rect 1448 103780 2147 103808
rect 2167 108162 2866 108190
rect 2167 103808 2782 108162
rect 2846 103808 2866 108162
rect 2167 103780 2866 103808
rect -2866 103652 -2167 103680
rect -2866 99298 -2251 103652
rect -2187 99298 -2167 103652
rect -2866 99270 -2167 99298
rect -2147 103652 -1448 103680
rect -2147 99298 -1532 103652
rect -1468 99298 -1448 103652
rect -2147 99270 -1448 99298
rect -1428 103652 -729 103680
rect -1428 99298 -813 103652
rect -749 99298 -729 103652
rect -1428 99270 -729 99298
rect -709 103652 -10 103680
rect -709 99298 -94 103652
rect -30 99298 -10 103652
rect -709 99270 -10 99298
rect 10 103652 709 103680
rect 10 99298 625 103652
rect 689 99298 709 103652
rect 10 99270 709 99298
rect 729 103652 1428 103680
rect 729 99298 1344 103652
rect 1408 99298 1428 103652
rect 729 99270 1428 99298
rect 1448 103652 2147 103680
rect 1448 99298 2063 103652
rect 2127 99298 2147 103652
rect 1448 99270 2147 99298
rect 2167 103652 2866 103680
rect 2167 99298 2782 103652
rect 2846 99298 2866 103652
rect 2167 99270 2866 99298
rect -2866 99142 -2167 99170
rect -2866 94788 -2251 99142
rect -2187 94788 -2167 99142
rect -2866 94760 -2167 94788
rect -2147 99142 -1448 99170
rect -2147 94788 -1532 99142
rect -1468 94788 -1448 99142
rect -2147 94760 -1448 94788
rect -1428 99142 -729 99170
rect -1428 94788 -813 99142
rect -749 94788 -729 99142
rect -1428 94760 -729 94788
rect -709 99142 -10 99170
rect -709 94788 -94 99142
rect -30 94788 -10 99142
rect -709 94760 -10 94788
rect 10 99142 709 99170
rect 10 94788 625 99142
rect 689 94788 709 99142
rect 10 94760 709 94788
rect 729 99142 1428 99170
rect 729 94788 1344 99142
rect 1408 94788 1428 99142
rect 729 94760 1428 94788
rect 1448 99142 2147 99170
rect 1448 94788 2063 99142
rect 2127 94788 2147 99142
rect 1448 94760 2147 94788
rect 2167 99142 2866 99170
rect 2167 94788 2782 99142
rect 2846 94788 2866 99142
rect 2167 94760 2866 94788
rect -2866 94632 -2167 94660
rect -2866 90278 -2251 94632
rect -2187 90278 -2167 94632
rect -2866 90250 -2167 90278
rect -2147 94632 -1448 94660
rect -2147 90278 -1532 94632
rect -1468 90278 -1448 94632
rect -2147 90250 -1448 90278
rect -1428 94632 -729 94660
rect -1428 90278 -813 94632
rect -749 90278 -729 94632
rect -1428 90250 -729 90278
rect -709 94632 -10 94660
rect -709 90278 -94 94632
rect -30 90278 -10 94632
rect -709 90250 -10 90278
rect 10 94632 709 94660
rect 10 90278 625 94632
rect 689 90278 709 94632
rect 10 90250 709 90278
rect 729 94632 1428 94660
rect 729 90278 1344 94632
rect 1408 90278 1428 94632
rect 729 90250 1428 90278
rect 1448 94632 2147 94660
rect 1448 90278 2063 94632
rect 2127 90278 2147 94632
rect 1448 90250 2147 90278
rect 2167 94632 2866 94660
rect 2167 90278 2782 94632
rect 2846 90278 2866 94632
rect 2167 90250 2866 90278
rect -2866 90122 -2167 90150
rect -2866 85768 -2251 90122
rect -2187 85768 -2167 90122
rect -2866 85740 -2167 85768
rect -2147 90122 -1448 90150
rect -2147 85768 -1532 90122
rect -1468 85768 -1448 90122
rect -2147 85740 -1448 85768
rect -1428 90122 -729 90150
rect -1428 85768 -813 90122
rect -749 85768 -729 90122
rect -1428 85740 -729 85768
rect -709 90122 -10 90150
rect -709 85768 -94 90122
rect -30 85768 -10 90122
rect -709 85740 -10 85768
rect 10 90122 709 90150
rect 10 85768 625 90122
rect 689 85768 709 90122
rect 10 85740 709 85768
rect 729 90122 1428 90150
rect 729 85768 1344 90122
rect 1408 85768 1428 90122
rect 729 85740 1428 85768
rect 1448 90122 2147 90150
rect 1448 85768 2063 90122
rect 2127 85768 2147 90122
rect 1448 85740 2147 85768
rect 2167 90122 2866 90150
rect 2167 85768 2782 90122
rect 2846 85768 2866 90122
rect 2167 85740 2866 85768
rect -2866 85612 -2167 85640
rect -2866 81258 -2251 85612
rect -2187 81258 -2167 85612
rect -2866 81230 -2167 81258
rect -2147 85612 -1448 85640
rect -2147 81258 -1532 85612
rect -1468 81258 -1448 85612
rect -2147 81230 -1448 81258
rect -1428 85612 -729 85640
rect -1428 81258 -813 85612
rect -749 81258 -729 85612
rect -1428 81230 -729 81258
rect -709 85612 -10 85640
rect -709 81258 -94 85612
rect -30 81258 -10 85612
rect -709 81230 -10 81258
rect 10 85612 709 85640
rect 10 81258 625 85612
rect 689 81258 709 85612
rect 10 81230 709 81258
rect 729 85612 1428 85640
rect 729 81258 1344 85612
rect 1408 81258 1428 85612
rect 729 81230 1428 81258
rect 1448 85612 2147 85640
rect 1448 81258 2063 85612
rect 2127 81258 2147 85612
rect 1448 81230 2147 81258
rect 2167 85612 2866 85640
rect 2167 81258 2782 85612
rect 2846 81258 2866 85612
rect 2167 81230 2866 81258
rect -2866 81102 -2167 81130
rect -2866 76748 -2251 81102
rect -2187 76748 -2167 81102
rect -2866 76720 -2167 76748
rect -2147 81102 -1448 81130
rect -2147 76748 -1532 81102
rect -1468 76748 -1448 81102
rect -2147 76720 -1448 76748
rect -1428 81102 -729 81130
rect -1428 76748 -813 81102
rect -749 76748 -729 81102
rect -1428 76720 -729 76748
rect -709 81102 -10 81130
rect -709 76748 -94 81102
rect -30 76748 -10 81102
rect -709 76720 -10 76748
rect 10 81102 709 81130
rect 10 76748 625 81102
rect 689 76748 709 81102
rect 10 76720 709 76748
rect 729 81102 1428 81130
rect 729 76748 1344 81102
rect 1408 76748 1428 81102
rect 729 76720 1428 76748
rect 1448 81102 2147 81130
rect 1448 76748 2063 81102
rect 2127 76748 2147 81102
rect 1448 76720 2147 76748
rect 2167 81102 2866 81130
rect 2167 76748 2782 81102
rect 2846 76748 2866 81102
rect 2167 76720 2866 76748
rect -2866 76592 -2167 76620
rect -2866 72238 -2251 76592
rect -2187 72238 -2167 76592
rect -2866 72210 -2167 72238
rect -2147 76592 -1448 76620
rect -2147 72238 -1532 76592
rect -1468 72238 -1448 76592
rect -2147 72210 -1448 72238
rect -1428 76592 -729 76620
rect -1428 72238 -813 76592
rect -749 72238 -729 76592
rect -1428 72210 -729 72238
rect -709 76592 -10 76620
rect -709 72238 -94 76592
rect -30 72238 -10 76592
rect -709 72210 -10 72238
rect 10 76592 709 76620
rect 10 72238 625 76592
rect 689 72238 709 76592
rect 10 72210 709 72238
rect 729 76592 1428 76620
rect 729 72238 1344 76592
rect 1408 72238 1428 76592
rect 729 72210 1428 72238
rect 1448 76592 2147 76620
rect 1448 72238 2063 76592
rect 2127 72238 2147 76592
rect 1448 72210 2147 72238
rect 2167 76592 2866 76620
rect 2167 72238 2782 76592
rect 2846 72238 2866 76592
rect 2167 72210 2866 72238
rect -2866 72082 -2167 72110
rect -2866 67728 -2251 72082
rect -2187 67728 -2167 72082
rect -2866 67700 -2167 67728
rect -2147 72082 -1448 72110
rect -2147 67728 -1532 72082
rect -1468 67728 -1448 72082
rect -2147 67700 -1448 67728
rect -1428 72082 -729 72110
rect -1428 67728 -813 72082
rect -749 67728 -729 72082
rect -1428 67700 -729 67728
rect -709 72082 -10 72110
rect -709 67728 -94 72082
rect -30 67728 -10 72082
rect -709 67700 -10 67728
rect 10 72082 709 72110
rect 10 67728 625 72082
rect 689 67728 709 72082
rect 10 67700 709 67728
rect 729 72082 1428 72110
rect 729 67728 1344 72082
rect 1408 67728 1428 72082
rect 729 67700 1428 67728
rect 1448 72082 2147 72110
rect 1448 67728 2063 72082
rect 2127 67728 2147 72082
rect 1448 67700 2147 67728
rect 2167 72082 2866 72110
rect 2167 67728 2782 72082
rect 2846 67728 2866 72082
rect 2167 67700 2866 67728
rect -2866 67572 -2167 67600
rect -2866 63218 -2251 67572
rect -2187 63218 -2167 67572
rect -2866 63190 -2167 63218
rect -2147 67572 -1448 67600
rect -2147 63218 -1532 67572
rect -1468 63218 -1448 67572
rect -2147 63190 -1448 63218
rect -1428 67572 -729 67600
rect -1428 63218 -813 67572
rect -749 63218 -729 67572
rect -1428 63190 -729 63218
rect -709 67572 -10 67600
rect -709 63218 -94 67572
rect -30 63218 -10 67572
rect -709 63190 -10 63218
rect 10 67572 709 67600
rect 10 63218 625 67572
rect 689 63218 709 67572
rect 10 63190 709 63218
rect 729 67572 1428 67600
rect 729 63218 1344 67572
rect 1408 63218 1428 67572
rect 729 63190 1428 63218
rect 1448 67572 2147 67600
rect 1448 63218 2063 67572
rect 2127 63218 2147 67572
rect 1448 63190 2147 63218
rect 2167 67572 2866 67600
rect 2167 63218 2782 67572
rect 2846 63218 2866 67572
rect 2167 63190 2866 63218
rect -2866 63062 -2167 63090
rect -2866 58708 -2251 63062
rect -2187 58708 -2167 63062
rect -2866 58680 -2167 58708
rect -2147 63062 -1448 63090
rect -2147 58708 -1532 63062
rect -1468 58708 -1448 63062
rect -2147 58680 -1448 58708
rect -1428 63062 -729 63090
rect -1428 58708 -813 63062
rect -749 58708 -729 63062
rect -1428 58680 -729 58708
rect -709 63062 -10 63090
rect -709 58708 -94 63062
rect -30 58708 -10 63062
rect -709 58680 -10 58708
rect 10 63062 709 63090
rect 10 58708 625 63062
rect 689 58708 709 63062
rect 10 58680 709 58708
rect 729 63062 1428 63090
rect 729 58708 1344 63062
rect 1408 58708 1428 63062
rect 729 58680 1428 58708
rect 1448 63062 2147 63090
rect 1448 58708 2063 63062
rect 2127 58708 2147 63062
rect 1448 58680 2147 58708
rect 2167 63062 2866 63090
rect 2167 58708 2782 63062
rect 2846 58708 2866 63062
rect 2167 58680 2866 58708
rect -2866 58552 -2167 58580
rect -2866 54198 -2251 58552
rect -2187 54198 -2167 58552
rect -2866 54170 -2167 54198
rect -2147 58552 -1448 58580
rect -2147 54198 -1532 58552
rect -1468 54198 -1448 58552
rect -2147 54170 -1448 54198
rect -1428 58552 -729 58580
rect -1428 54198 -813 58552
rect -749 54198 -729 58552
rect -1428 54170 -729 54198
rect -709 58552 -10 58580
rect -709 54198 -94 58552
rect -30 54198 -10 58552
rect -709 54170 -10 54198
rect 10 58552 709 58580
rect 10 54198 625 58552
rect 689 54198 709 58552
rect 10 54170 709 54198
rect 729 58552 1428 58580
rect 729 54198 1344 58552
rect 1408 54198 1428 58552
rect 729 54170 1428 54198
rect 1448 58552 2147 58580
rect 1448 54198 2063 58552
rect 2127 54198 2147 58552
rect 1448 54170 2147 54198
rect 2167 58552 2866 58580
rect 2167 54198 2782 58552
rect 2846 54198 2866 58552
rect 2167 54170 2866 54198
rect -2866 54042 -2167 54070
rect -2866 49688 -2251 54042
rect -2187 49688 -2167 54042
rect -2866 49660 -2167 49688
rect -2147 54042 -1448 54070
rect -2147 49688 -1532 54042
rect -1468 49688 -1448 54042
rect -2147 49660 -1448 49688
rect -1428 54042 -729 54070
rect -1428 49688 -813 54042
rect -749 49688 -729 54042
rect -1428 49660 -729 49688
rect -709 54042 -10 54070
rect -709 49688 -94 54042
rect -30 49688 -10 54042
rect -709 49660 -10 49688
rect 10 54042 709 54070
rect 10 49688 625 54042
rect 689 49688 709 54042
rect 10 49660 709 49688
rect 729 54042 1428 54070
rect 729 49688 1344 54042
rect 1408 49688 1428 54042
rect 729 49660 1428 49688
rect 1448 54042 2147 54070
rect 1448 49688 2063 54042
rect 2127 49688 2147 54042
rect 1448 49660 2147 49688
rect 2167 54042 2866 54070
rect 2167 49688 2782 54042
rect 2846 49688 2866 54042
rect 2167 49660 2866 49688
rect -2866 49532 -2167 49560
rect -2866 45178 -2251 49532
rect -2187 45178 -2167 49532
rect -2866 45150 -2167 45178
rect -2147 49532 -1448 49560
rect -2147 45178 -1532 49532
rect -1468 45178 -1448 49532
rect -2147 45150 -1448 45178
rect -1428 49532 -729 49560
rect -1428 45178 -813 49532
rect -749 45178 -729 49532
rect -1428 45150 -729 45178
rect -709 49532 -10 49560
rect -709 45178 -94 49532
rect -30 45178 -10 49532
rect -709 45150 -10 45178
rect 10 49532 709 49560
rect 10 45178 625 49532
rect 689 45178 709 49532
rect 10 45150 709 45178
rect 729 49532 1428 49560
rect 729 45178 1344 49532
rect 1408 45178 1428 49532
rect 729 45150 1428 45178
rect 1448 49532 2147 49560
rect 1448 45178 2063 49532
rect 2127 45178 2147 49532
rect 1448 45150 2147 45178
rect 2167 49532 2866 49560
rect 2167 45178 2782 49532
rect 2846 45178 2866 49532
rect 2167 45150 2866 45178
rect -2866 45022 -2167 45050
rect -2866 40668 -2251 45022
rect -2187 40668 -2167 45022
rect -2866 40640 -2167 40668
rect -2147 45022 -1448 45050
rect -2147 40668 -1532 45022
rect -1468 40668 -1448 45022
rect -2147 40640 -1448 40668
rect -1428 45022 -729 45050
rect -1428 40668 -813 45022
rect -749 40668 -729 45022
rect -1428 40640 -729 40668
rect -709 45022 -10 45050
rect -709 40668 -94 45022
rect -30 40668 -10 45022
rect -709 40640 -10 40668
rect 10 45022 709 45050
rect 10 40668 625 45022
rect 689 40668 709 45022
rect 10 40640 709 40668
rect 729 45022 1428 45050
rect 729 40668 1344 45022
rect 1408 40668 1428 45022
rect 729 40640 1428 40668
rect 1448 45022 2147 45050
rect 1448 40668 2063 45022
rect 2127 40668 2147 45022
rect 1448 40640 2147 40668
rect 2167 45022 2866 45050
rect 2167 40668 2782 45022
rect 2846 40668 2866 45022
rect 2167 40640 2866 40668
rect -2866 40512 -2167 40540
rect -2866 36158 -2251 40512
rect -2187 36158 -2167 40512
rect -2866 36130 -2167 36158
rect -2147 40512 -1448 40540
rect -2147 36158 -1532 40512
rect -1468 36158 -1448 40512
rect -2147 36130 -1448 36158
rect -1428 40512 -729 40540
rect -1428 36158 -813 40512
rect -749 36158 -729 40512
rect -1428 36130 -729 36158
rect -709 40512 -10 40540
rect -709 36158 -94 40512
rect -30 36158 -10 40512
rect -709 36130 -10 36158
rect 10 40512 709 40540
rect 10 36158 625 40512
rect 689 36158 709 40512
rect 10 36130 709 36158
rect 729 40512 1428 40540
rect 729 36158 1344 40512
rect 1408 36158 1428 40512
rect 729 36130 1428 36158
rect 1448 40512 2147 40540
rect 1448 36158 2063 40512
rect 2127 36158 2147 40512
rect 1448 36130 2147 36158
rect 2167 40512 2866 40540
rect 2167 36158 2782 40512
rect 2846 36158 2866 40512
rect 2167 36130 2866 36158
rect -2866 36002 -2167 36030
rect -2866 31648 -2251 36002
rect -2187 31648 -2167 36002
rect -2866 31620 -2167 31648
rect -2147 36002 -1448 36030
rect -2147 31648 -1532 36002
rect -1468 31648 -1448 36002
rect -2147 31620 -1448 31648
rect -1428 36002 -729 36030
rect -1428 31648 -813 36002
rect -749 31648 -729 36002
rect -1428 31620 -729 31648
rect -709 36002 -10 36030
rect -709 31648 -94 36002
rect -30 31648 -10 36002
rect -709 31620 -10 31648
rect 10 36002 709 36030
rect 10 31648 625 36002
rect 689 31648 709 36002
rect 10 31620 709 31648
rect 729 36002 1428 36030
rect 729 31648 1344 36002
rect 1408 31648 1428 36002
rect 729 31620 1428 31648
rect 1448 36002 2147 36030
rect 1448 31648 2063 36002
rect 2127 31648 2147 36002
rect 1448 31620 2147 31648
rect 2167 36002 2866 36030
rect 2167 31648 2782 36002
rect 2846 31648 2866 36002
rect 2167 31620 2866 31648
rect -2866 31492 -2167 31520
rect -2866 27138 -2251 31492
rect -2187 27138 -2167 31492
rect -2866 27110 -2167 27138
rect -2147 31492 -1448 31520
rect -2147 27138 -1532 31492
rect -1468 27138 -1448 31492
rect -2147 27110 -1448 27138
rect -1428 31492 -729 31520
rect -1428 27138 -813 31492
rect -749 27138 -729 31492
rect -1428 27110 -729 27138
rect -709 31492 -10 31520
rect -709 27138 -94 31492
rect -30 27138 -10 31492
rect -709 27110 -10 27138
rect 10 31492 709 31520
rect 10 27138 625 31492
rect 689 27138 709 31492
rect 10 27110 709 27138
rect 729 31492 1428 31520
rect 729 27138 1344 31492
rect 1408 27138 1428 31492
rect 729 27110 1428 27138
rect 1448 31492 2147 31520
rect 1448 27138 2063 31492
rect 2127 27138 2147 31492
rect 1448 27110 2147 27138
rect 2167 31492 2866 31520
rect 2167 27138 2782 31492
rect 2846 27138 2866 31492
rect 2167 27110 2866 27138
rect -2866 26982 -2167 27010
rect -2866 22628 -2251 26982
rect -2187 22628 -2167 26982
rect -2866 22600 -2167 22628
rect -2147 26982 -1448 27010
rect -2147 22628 -1532 26982
rect -1468 22628 -1448 26982
rect -2147 22600 -1448 22628
rect -1428 26982 -729 27010
rect -1428 22628 -813 26982
rect -749 22628 -729 26982
rect -1428 22600 -729 22628
rect -709 26982 -10 27010
rect -709 22628 -94 26982
rect -30 22628 -10 26982
rect -709 22600 -10 22628
rect 10 26982 709 27010
rect 10 22628 625 26982
rect 689 22628 709 26982
rect 10 22600 709 22628
rect 729 26982 1428 27010
rect 729 22628 1344 26982
rect 1408 22628 1428 26982
rect 729 22600 1428 22628
rect 1448 26982 2147 27010
rect 1448 22628 2063 26982
rect 2127 22628 2147 26982
rect 1448 22600 2147 22628
rect 2167 26982 2866 27010
rect 2167 22628 2782 26982
rect 2846 22628 2866 26982
rect 2167 22600 2866 22628
rect -2866 22472 -2167 22500
rect -2866 18118 -2251 22472
rect -2187 18118 -2167 22472
rect -2866 18090 -2167 18118
rect -2147 22472 -1448 22500
rect -2147 18118 -1532 22472
rect -1468 18118 -1448 22472
rect -2147 18090 -1448 18118
rect -1428 22472 -729 22500
rect -1428 18118 -813 22472
rect -749 18118 -729 22472
rect -1428 18090 -729 18118
rect -709 22472 -10 22500
rect -709 18118 -94 22472
rect -30 18118 -10 22472
rect -709 18090 -10 18118
rect 10 22472 709 22500
rect 10 18118 625 22472
rect 689 18118 709 22472
rect 10 18090 709 18118
rect 729 22472 1428 22500
rect 729 18118 1344 22472
rect 1408 18118 1428 22472
rect 729 18090 1428 18118
rect 1448 22472 2147 22500
rect 1448 18118 2063 22472
rect 2127 18118 2147 22472
rect 1448 18090 2147 18118
rect 2167 22472 2866 22500
rect 2167 18118 2782 22472
rect 2846 18118 2866 22472
rect 2167 18090 2866 18118
rect -2866 17962 -2167 17990
rect -2866 13608 -2251 17962
rect -2187 13608 -2167 17962
rect -2866 13580 -2167 13608
rect -2147 17962 -1448 17990
rect -2147 13608 -1532 17962
rect -1468 13608 -1448 17962
rect -2147 13580 -1448 13608
rect -1428 17962 -729 17990
rect -1428 13608 -813 17962
rect -749 13608 -729 17962
rect -1428 13580 -729 13608
rect -709 17962 -10 17990
rect -709 13608 -94 17962
rect -30 13608 -10 17962
rect -709 13580 -10 13608
rect 10 17962 709 17990
rect 10 13608 625 17962
rect 689 13608 709 17962
rect 10 13580 709 13608
rect 729 17962 1428 17990
rect 729 13608 1344 17962
rect 1408 13608 1428 17962
rect 729 13580 1428 13608
rect 1448 17962 2147 17990
rect 1448 13608 2063 17962
rect 2127 13608 2147 17962
rect 1448 13580 2147 13608
rect 2167 17962 2866 17990
rect 2167 13608 2782 17962
rect 2846 13608 2866 17962
rect 2167 13580 2866 13608
rect -2866 13452 -2167 13480
rect -2866 9098 -2251 13452
rect -2187 9098 -2167 13452
rect -2866 9070 -2167 9098
rect -2147 13452 -1448 13480
rect -2147 9098 -1532 13452
rect -1468 9098 -1448 13452
rect -2147 9070 -1448 9098
rect -1428 13452 -729 13480
rect -1428 9098 -813 13452
rect -749 9098 -729 13452
rect -1428 9070 -729 9098
rect -709 13452 -10 13480
rect -709 9098 -94 13452
rect -30 9098 -10 13452
rect -709 9070 -10 9098
rect 10 13452 709 13480
rect 10 9098 625 13452
rect 689 9098 709 13452
rect 10 9070 709 9098
rect 729 13452 1428 13480
rect 729 9098 1344 13452
rect 1408 9098 1428 13452
rect 729 9070 1428 9098
rect 1448 13452 2147 13480
rect 1448 9098 2063 13452
rect 2127 9098 2147 13452
rect 1448 9070 2147 9098
rect 2167 13452 2866 13480
rect 2167 9098 2782 13452
rect 2846 9098 2866 13452
rect 2167 9070 2866 9098
rect -2866 8942 -2167 8970
rect -2866 4588 -2251 8942
rect -2187 4588 -2167 8942
rect -2866 4560 -2167 4588
rect -2147 8942 -1448 8970
rect -2147 4588 -1532 8942
rect -1468 4588 -1448 8942
rect -2147 4560 -1448 4588
rect -1428 8942 -729 8970
rect -1428 4588 -813 8942
rect -749 4588 -729 8942
rect -1428 4560 -729 4588
rect -709 8942 -10 8970
rect -709 4588 -94 8942
rect -30 4588 -10 8942
rect -709 4560 -10 4588
rect 10 8942 709 8970
rect 10 4588 625 8942
rect 689 4588 709 8942
rect 10 4560 709 4588
rect 729 8942 1428 8970
rect 729 4588 1344 8942
rect 1408 4588 1428 8942
rect 729 4560 1428 4588
rect 1448 8942 2147 8970
rect 1448 4588 2063 8942
rect 2127 4588 2147 8942
rect 1448 4560 2147 4588
rect 2167 8942 2866 8970
rect 2167 4588 2782 8942
rect 2846 4588 2866 8942
rect 2167 4560 2866 4588
rect -2866 4432 -2167 4460
rect -2866 78 -2251 4432
rect -2187 78 -2167 4432
rect -2866 50 -2167 78
rect -2147 4432 -1448 4460
rect -2147 78 -1532 4432
rect -1468 78 -1448 4432
rect -2147 50 -1448 78
rect -1428 4432 -729 4460
rect -1428 78 -813 4432
rect -749 78 -729 4432
rect -1428 50 -729 78
rect -709 4432 -10 4460
rect -709 78 -94 4432
rect -30 78 -10 4432
rect -709 50 -10 78
rect 10 4432 709 4460
rect 10 78 625 4432
rect 689 78 709 4432
rect 10 50 709 78
rect 729 4432 1428 4460
rect 729 78 1344 4432
rect 1408 78 1428 4432
rect 729 50 1428 78
rect 1448 4432 2147 4460
rect 1448 78 2063 4432
rect 2127 78 2147 4432
rect 1448 50 2147 78
rect 2167 4432 2866 4460
rect 2167 78 2782 4432
rect 2846 78 2866 4432
rect 2167 50 2866 78
rect -2866 -78 -2167 -50
rect -2866 -4432 -2251 -78
rect -2187 -4432 -2167 -78
rect -2866 -4460 -2167 -4432
rect -2147 -78 -1448 -50
rect -2147 -4432 -1532 -78
rect -1468 -4432 -1448 -78
rect -2147 -4460 -1448 -4432
rect -1428 -78 -729 -50
rect -1428 -4432 -813 -78
rect -749 -4432 -729 -78
rect -1428 -4460 -729 -4432
rect -709 -78 -10 -50
rect -709 -4432 -94 -78
rect -30 -4432 -10 -78
rect -709 -4460 -10 -4432
rect 10 -78 709 -50
rect 10 -4432 625 -78
rect 689 -4432 709 -78
rect 10 -4460 709 -4432
rect 729 -78 1428 -50
rect 729 -4432 1344 -78
rect 1408 -4432 1428 -78
rect 729 -4460 1428 -4432
rect 1448 -78 2147 -50
rect 1448 -4432 2063 -78
rect 2127 -4432 2147 -78
rect 1448 -4460 2147 -4432
rect 2167 -78 2866 -50
rect 2167 -4432 2782 -78
rect 2846 -4432 2866 -78
rect 2167 -4460 2866 -4432
rect -2866 -4588 -2167 -4560
rect -2866 -8942 -2251 -4588
rect -2187 -8942 -2167 -4588
rect -2866 -8970 -2167 -8942
rect -2147 -4588 -1448 -4560
rect -2147 -8942 -1532 -4588
rect -1468 -8942 -1448 -4588
rect -2147 -8970 -1448 -8942
rect -1428 -4588 -729 -4560
rect -1428 -8942 -813 -4588
rect -749 -8942 -729 -4588
rect -1428 -8970 -729 -8942
rect -709 -4588 -10 -4560
rect -709 -8942 -94 -4588
rect -30 -8942 -10 -4588
rect -709 -8970 -10 -8942
rect 10 -4588 709 -4560
rect 10 -8942 625 -4588
rect 689 -8942 709 -4588
rect 10 -8970 709 -8942
rect 729 -4588 1428 -4560
rect 729 -8942 1344 -4588
rect 1408 -8942 1428 -4588
rect 729 -8970 1428 -8942
rect 1448 -4588 2147 -4560
rect 1448 -8942 2063 -4588
rect 2127 -8942 2147 -4588
rect 1448 -8970 2147 -8942
rect 2167 -4588 2866 -4560
rect 2167 -8942 2782 -4588
rect 2846 -8942 2866 -4588
rect 2167 -8970 2866 -8942
rect -2866 -9098 -2167 -9070
rect -2866 -13452 -2251 -9098
rect -2187 -13452 -2167 -9098
rect -2866 -13480 -2167 -13452
rect -2147 -9098 -1448 -9070
rect -2147 -13452 -1532 -9098
rect -1468 -13452 -1448 -9098
rect -2147 -13480 -1448 -13452
rect -1428 -9098 -729 -9070
rect -1428 -13452 -813 -9098
rect -749 -13452 -729 -9098
rect -1428 -13480 -729 -13452
rect -709 -9098 -10 -9070
rect -709 -13452 -94 -9098
rect -30 -13452 -10 -9098
rect -709 -13480 -10 -13452
rect 10 -9098 709 -9070
rect 10 -13452 625 -9098
rect 689 -13452 709 -9098
rect 10 -13480 709 -13452
rect 729 -9098 1428 -9070
rect 729 -13452 1344 -9098
rect 1408 -13452 1428 -9098
rect 729 -13480 1428 -13452
rect 1448 -9098 2147 -9070
rect 1448 -13452 2063 -9098
rect 2127 -13452 2147 -9098
rect 1448 -13480 2147 -13452
rect 2167 -9098 2866 -9070
rect 2167 -13452 2782 -9098
rect 2846 -13452 2866 -9098
rect 2167 -13480 2866 -13452
rect -2866 -13608 -2167 -13580
rect -2866 -17962 -2251 -13608
rect -2187 -17962 -2167 -13608
rect -2866 -17990 -2167 -17962
rect -2147 -13608 -1448 -13580
rect -2147 -17962 -1532 -13608
rect -1468 -17962 -1448 -13608
rect -2147 -17990 -1448 -17962
rect -1428 -13608 -729 -13580
rect -1428 -17962 -813 -13608
rect -749 -17962 -729 -13608
rect -1428 -17990 -729 -17962
rect -709 -13608 -10 -13580
rect -709 -17962 -94 -13608
rect -30 -17962 -10 -13608
rect -709 -17990 -10 -17962
rect 10 -13608 709 -13580
rect 10 -17962 625 -13608
rect 689 -17962 709 -13608
rect 10 -17990 709 -17962
rect 729 -13608 1428 -13580
rect 729 -17962 1344 -13608
rect 1408 -17962 1428 -13608
rect 729 -17990 1428 -17962
rect 1448 -13608 2147 -13580
rect 1448 -17962 2063 -13608
rect 2127 -17962 2147 -13608
rect 1448 -17990 2147 -17962
rect 2167 -13608 2866 -13580
rect 2167 -17962 2782 -13608
rect 2846 -17962 2866 -13608
rect 2167 -17990 2866 -17962
rect -2866 -18118 -2167 -18090
rect -2866 -22472 -2251 -18118
rect -2187 -22472 -2167 -18118
rect -2866 -22500 -2167 -22472
rect -2147 -18118 -1448 -18090
rect -2147 -22472 -1532 -18118
rect -1468 -22472 -1448 -18118
rect -2147 -22500 -1448 -22472
rect -1428 -18118 -729 -18090
rect -1428 -22472 -813 -18118
rect -749 -22472 -729 -18118
rect -1428 -22500 -729 -22472
rect -709 -18118 -10 -18090
rect -709 -22472 -94 -18118
rect -30 -22472 -10 -18118
rect -709 -22500 -10 -22472
rect 10 -18118 709 -18090
rect 10 -22472 625 -18118
rect 689 -22472 709 -18118
rect 10 -22500 709 -22472
rect 729 -18118 1428 -18090
rect 729 -22472 1344 -18118
rect 1408 -22472 1428 -18118
rect 729 -22500 1428 -22472
rect 1448 -18118 2147 -18090
rect 1448 -22472 2063 -18118
rect 2127 -22472 2147 -18118
rect 1448 -22500 2147 -22472
rect 2167 -18118 2866 -18090
rect 2167 -22472 2782 -18118
rect 2846 -22472 2866 -18118
rect 2167 -22500 2866 -22472
rect -2866 -22628 -2167 -22600
rect -2866 -26982 -2251 -22628
rect -2187 -26982 -2167 -22628
rect -2866 -27010 -2167 -26982
rect -2147 -22628 -1448 -22600
rect -2147 -26982 -1532 -22628
rect -1468 -26982 -1448 -22628
rect -2147 -27010 -1448 -26982
rect -1428 -22628 -729 -22600
rect -1428 -26982 -813 -22628
rect -749 -26982 -729 -22628
rect -1428 -27010 -729 -26982
rect -709 -22628 -10 -22600
rect -709 -26982 -94 -22628
rect -30 -26982 -10 -22628
rect -709 -27010 -10 -26982
rect 10 -22628 709 -22600
rect 10 -26982 625 -22628
rect 689 -26982 709 -22628
rect 10 -27010 709 -26982
rect 729 -22628 1428 -22600
rect 729 -26982 1344 -22628
rect 1408 -26982 1428 -22628
rect 729 -27010 1428 -26982
rect 1448 -22628 2147 -22600
rect 1448 -26982 2063 -22628
rect 2127 -26982 2147 -22628
rect 1448 -27010 2147 -26982
rect 2167 -22628 2866 -22600
rect 2167 -26982 2782 -22628
rect 2846 -26982 2866 -22628
rect 2167 -27010 2866 -26982
rect -2866 -27138 -2167 -27110
rect -2866 -31492 -2251 -27138
rect -2187 -31492 -2167 -27138
rect -2866 -31520 -2167 -31492
rect -2147 -27138 -1448 -27110
rect -2147 -31492 -1532 -27138
rect -1468 -31492 -1448 -27138
rect -2147 -31520 -1448 -31492
rect -1428 -27138 -729 -27110
rect -1428 -31492 -813 -27138
rect -749 -31492 -729 -27138
rect -1428 -31520 -729 -31492
rect -709 -27138 -10 -27110
rect -709 -31492 -94 -27138
rect -30 -31492 -10 -27138
rect -709 -31520 -10 -31492
rect 10 -27138 709 -27110
rect 10 -31492 625 -27138
rect 689 -31492 709 -27138
rect 10 -31520 709 -31492
rect 729 -27138 1428 -27110
rect 729 -31492 1344 -27138
rect 1408 -31492 1428 -27138
rect 729 -31520 1428 -31492
rect 1448 -27138 2147 -27110
rect 1448 -31492 2063 -27138
rect 2127 -31492 2147 -27138
rect 1448 -31520 2147 -31492
rect 2167 -27138 2866 -27110
rect 2167 -31492 2782 -27138
rect 2846 -31492 2866 -27138
rect 2167 -31520 2866 -31492
rect -2866 -31648 -2167 -31620
rect -2866 -36002 -2251 -31648
rect -2187 -36002 -2167 -31648
rect -2866 -36030 -2167 -36002
rect -2147 -31648 -1448 -31620
rect -2147 -36002 -1532 -31648
rect -1468 -36002 -1448 -31648
rect -2147 -36030 -1448 -36002
rect -1428 -31648 -729 -31620
rect -1428 -36002 -813 -31648
rect -749 -36002 -729 -31648
rect -1428 -36030 -729 -36002
rect -709 -31648 -10 -31620
rect -709 -36002 -94 -31648
rect -30 -36002 -10 -31648
rect -709 -36030 -10 -36002
rect 10 -31648 709 -31620
rect 10 -36002 625 -31648
rect 689 -36002 709 -31648
rect 10 -36030 709 -36002
rect 729 -31648 1428 -31620
rect 729 -36002 1344 -31648
rect 1408 -36002 1428 -31648
rect 729 -36030 1428 -36002
rect 1448 -31648 2147 -31620
rect 1448 -36002 2063 -31648
rect 2127 -36002 2147 -31648
rect 1448 -36030 2147 -36002
rect 2167 -31648 2866 -31620
rect 2167 -36002 2782 -31648
rect 2846 -36002 2866 -31648
rect 2167 -36030 2866 -36002
rect -2866 -36158 -2167 -36130
rect -2866 -40512 -2251 -36158
rect -2187 -40512 -2167 -36158
rect -2866 -40540 -2167 -40512
rect -2147 -36158 -1448 -36130
rect -2147 -40512 -1532 -36158
rect -1468 -40512 -1448 -36158
rect -2147 -40540 -1448 -40512
rect -1428 -36158 -729 -36130
rect -1428 -40512 -813 -36158
rect -749 -40512 -729 -36158
rect -1428 -40540 -729 -40512
rect -709 -36158 -10 -36130
rect -709 -40512 -94 -36158
rect -30 -40512 -10 -36158
rect -709 -40540 -10 -40512
rect 10 -36158 709 -36130
rect 10 -40512 625 -36158
rect 689 -40512 709 -36158
rect 10 -40540 709 -40512
rect 729 -36158 1428 -36130
rect 729 -40512 1344 -36158
rect 1408 -40512 1428 -36158
rect 729 -40540 1428 -40512
rect 1448 -36158 2147 -36130
rect 1448 -40512 2063 -36158
rect 2127 -40512 2147 -36158
rect 1448 -40540 2147 -40512
rect 2167 -36158 2866 -36130
rect 2167 -40512 2782 -36158
rect 2846 -40512 2866 -36158
rect 2167 -40540 2866 -40512
rect -2866 -40668 -2167 -40640
rect -2866 -45022 -2251 -40668
rect -2187 -45022 -2167 -40668
rect -2866 -45050 -2167 -45022
rect -2147 -40668 -1448 -40640
rect -2147 -45022 -1532 -40668
rect -1468 -45022 -1448 -40668
rect -2147 -45050 -1448 -45022
rect -1428 -40668 -729 -40640
rect -1428 -45022 -813 -40668
rect -749 -45022 -729 -40668
rect -1428 -45050 -729 -45022
rect -709 -40668 -10 -40640
rect -709 -45022 -94 -40668
rect -30 -45022 -10 -40668
rect -709 -45050 -10 -45022
rect 10 -40668 709 -40640
rect 10 -45022 625 -40668
rect 689 -45022 709 -40668
rect 10 -45050 709 -45022
rect 729 -40668 1428 -40640
rect 729 -45022 1344 -40668
rect 1408 -45022 1428 -40668
rect 729 -45050 1428 -45022
rect 1448 -40668 2147 -40640
rect 1448 -45022 2063 -40668
rect 2127 -45022 2147 -40668
rect 1448 -45050 2147 -45022
rect 2167 -40668 2866 -40640
rect 2167 -45022 2782 -40668
rect 2846 -45022 2866 -40668
rect 2167 -45050 2866 -45022
rect -2866 -45178 -2167 -45150
rect -2866 -49532 -2251 -45178
rect -2187 -49532 -2167 -45178
rect -2866 -49560 -2167 -49532
rect -2147 -45178 -1448 -45150
rect -2147 -49532 -1532 -45178
rect -1468 -49532 -1448 -45178
rect -2147 -49560 -1448 -49532
rect -1428 -45178 -729 -45150
rect -1428 -49532 -813 -45178
rect -749 -49532 -729 -45178
rect -1428 -49560 -729 -49532
rect -709 -45178 -10 -45150
rect -709 -49532 -94 -45178
rect -30 -49532 -10 -45178
rect -709 -49560 -10 -49532
rect 10 -45178 709 -45150
rect 10 -49532 625 -45178
rect 689 -49532 709 -45178
rect 10 -49560 709 -49532
rect 729 -45178 1428 -45150
rect 729 -49532 1344 -45178
rect 1408 -49532 1428 -45178
rect 729 -49560 1428 -49532
rect 1448 -45178 2147 -45150
rect 1448 -49532 2063 -45178
rect 2127 -49532 2147 -45178
rect 1448 -49560 2147 -49532
rect 2167 -45178 2866 -45150
rect 2167 -49532 2782 -45178
rect 2846 -49532 2866 -45178
rect 2167 -49560 2866 -49532
rect -2866 -49688 -2167 -49660
rect -2866 -54042 -2251 -49688
rect -2187 -54042 -2167 -49688
rect -2866 -54070 -2167 -54042
rect -2147 -49688 -1448 -49660
rect -2147 -54042 -1532 -49688
rect -1468 -54042 -1448 -49688
rect -2147 -54070 -1448 -54042
rect -1428 -49688 -729 -49660
rect -1428 -54042 -813 -49688
rect -749 -54042 -729 -49688
rect -1428 -54070 -729 -54042
rect -709 -49688 -10 -49660
rect -709 -54042 -94 -49688
rect -30 -54042 -10 -49688
rect -709 -54070 -10 -54042
rect 10 -49688 709 -49660
rect 10 -54042 625 -49688
rect 689 -54042 709 -49688
rect 10 -54070 709 -54042
rect 729 -49688 1428 -49660
rect 729 -54042 1344 -49688
rect 1408 -54042 1428 -49688
rect 729 -54070 1428 -54042
rect 1448 -49688 2147 -49660
rect 1448 -54042 2063 -49688
rect 2127 -54042 2147 -49688
rect 1448 -54070 2147 -54042
rect 2167 -49688 2866 -49660
rect 2167 -54042 2782 -49688
rect 2846 -54042 2866 -49688
rect 2167 -54070 2866 -54042
rect -2866 -54198 -2167 -54170
rect -2866 -58552 -2251 -54198
rect -2187 -58552 -2167 -54198
rect -2866 -58580 -2167 -58552
rect -2147 -54198 -1448 -54170
rect -2147 -58552 -1532 -54198
rect -1468 -58552 -1448 -54198
rect -2147 -58580 -1448 -58552
rect -1428 -54198 -729 -54170
rect -1428 -58552 -813 -54198
rect -749 -58552 -729 -54198
rect -1428 -58580 -729 -58552
rect -709 -54198 -10 -54170
rect -709 -58552 -94 -54198
rect -30 -58552 -10 -54198
rect -709 -58580 -10 -58552
rect 10 -54198 709 -54170
rect 10 -58552 625 -54198
rect 689 -58552 709 -54198
rect 10 -58580 709 -58552
rect 729 -54198 1428 -54170
rect 729 -58552 1344 -54198
rect 1408 -58552 1428 -54198
rect 729 -58580 1428 -58552
rect 1448 -54198 2147 -54170
rect 1448 -58552 2063 -54198
rect 2127 -58552 2147 -54198
rect 1448 -58580 2147 -58552
rect 2167 -54198 2866 -54170
rect 2167 -58552 2782 -54198
rect 2846 -58552 2866 -54198
rect 2167 -58580 2866 -58552
rect -2866 -58708 -2167 -58680
rect -2866 -63062 -2251 -58708
rect -2187 -63062 -2167 -58708
rect -2866 -63090 -2167 -63062
rect -2147 -58708 -1448 -58680
rect -2147 -63062 -1532 -58708
rect -1468 -63062 -1448 -58708
rect -2147 -63090 -1448 -63062
rect -1428 -58708 -729 -58680
rect -1428 -63062 -813 -58708
rect -749 -63062 -729 -58708
rect -1428 -63090 -729 -63062
rect -709 -58708 -10 -58680
rect -709 -63062 -94 -58708
rect -30 -63062 -10 -58708
rect -709 -63090 -10 -63062
rect 10 -58708 709 -58680
rect 10 -63062 625 -58708
rect 689 -63062 709 -58708
rect 10 -63090 709 -63062
rect 729 -58708 1428 -58680
rect 729 -63062 1344 -58708
rect 1408 -63062 1428 -58708
rect 729 -63090 1428 -63062
rect 1448 -58708 2147 -58680
rect 1448 -63062 2063 -58708
rect 2127 -63062 2147 -58708
rect 1448 -63090 2147 -63062
rect 2167 -58708 2866 -58680
rect 2167 -63062 2782 -58708
rect 2846 -63062 2866 -58708
rect 2167 -63090 2866 -63062
rect -2866 -63218 -2167 -63190
rect -2866 -67572 -2251 -63218
rect -2187 -67572 -2167 -63218
rect -2866 -67600 -2167 -67572
rect -2147 -63218 -1448 -63190
rect -2147 -67572 -1532 -63218
rect -1468 -67572 -1448 -63218
rect -2147 -67600 -1448 -67572
rect -1428 -63218 -729 -63190
rect -1428 -67572 -813 -63218
rect -749 -67572 -729 -63218
rect -1428 -67600 -729 -67572
rect -709 -63218 -10 -63190
rect -709 -67572 -94 -63218
rect -30 -67572 -10 -63218
rect -709 -67600 -10 -67572
rect 10 -63218 709 -63190
rect 10 -67572 625 -63218
rect 689 -67572 709 -63218
rect 10 -67600 709 -67572
rect 729 -63218 1428 -63190
rect 729 -67572 1344 -63218
rect 1408 -67572 1428 -63218
rect 729 -67600 1428 -67572
rect 1448 -63218 2147 -63190
rect 1448 -67572 2063 -63218
rect 2127 -67572 2147 -63218
rect 1448 -67600 2147 -67572
rect 2167 -63218 2866 -63190
rect 2167 -67572 2782 -63218
rect 2846 -67572 2866 -63218
rect 2167 -67600 2866 -67572
rect -2866 -67728 -2167 -67700
rect -2866 -72082 -2251 -67728
rect -2187 -72082 -2167 -67728
rect -2866 -72110 -2167 -72082
rect -2147 -67728 -1448 -67700
rect -2147 -72082 -1532 -67728
rect -1468 -72082 -1448 -67728
rect -2147 -72110 -1448 -72082
rect -1428 -67728 -729 -67700
rect -1428 -72082 -813 -67728
rect -749 -72082 -729 -67728
rect -1428 -72110 -729 -72082
rect -709 -67728 -10 -67700
rect -709 -72082 -94 -67728
rect -30 -72082 -10 -67728
rect -709 -72110 -10 -72082
rect 10 -67728 709 -67700
rect 10 -72082 625 -67728
rect 689 -72082 709 -67728
rect 10 -72110 709 -72082
rect 729 -67728 1428 -67700
rect 729 -72082 1344 -67728
rect 1408 -72082 1428 -67728
rect 729 -72110 1428 -72082
rect 1448 -67728 2147 -67700
rect 1448 -72082 2063 -67728
rect 2127 -72082 2147 -67728
rect 1448 -72110 2147 -72082
rect 2167 -67728 2866 -67700
rect 2167 -72082 2782 -67728
rect 2846 -72082 2866 -67728
rect 2167 -72110 2866 -72082
rect -2866 -72238 -2167 -72210
rect -2866 -76592 -2251 -72238
rect -2187 -76592 -2167 -72238
rect -2866 -76620 -2167 -76592
rect -2147 -72238 -1448 -72210
rect -2147 -76592 -1532 -72238
rect -1468 -76592 -1448 -72238
rect -2147 -76620 -1448 -76592
rect -1428 -72238 -729 -72210
rect -1428 -76592 -813 -72238
rect -749 -76592 -729 -72238
rect -1428 -76620 -729 -76592
rect -709 -72238 -10 -72210
rect -709 -76592 -94 -72238
rect -30 -76592 -10 -72238
rect -709 -76620 -10 -76592
rect 10 -72238 709 -72210
rect 10 -76592 625 -72238
rect 689 -76592 709 -72238
rect 10 -76620 709 -76592
rect 729 -72238 1428 -72210
rect 729 -76592 1344 -72238
rect 1408 -76592 1428 -72238
rect 729 -76620 1428 -76592
rect 1448 -72238 2147 -72210
rect 1448 -76592 2063 -72238
rect 2127 -76592 2147 -72238
rect 1448 -76620 2147 -76592
rect 2167 -72238 2866 -72210
rect 2167 -76592 2782 -72238
rect 2846 -76592 2866 -72238
rect 2167 -76620 2866 -76592
rect -2866 -76748 -2167 -76720
rect -2866 -81102 -2251 -76748
rect -2187 -81102 -2167 -76748
rect -2866 -81130 -2167 -81102
rect -2147 -76748 -1448 -76720
rect -2147 -81102 -1532 -76748
rect -1468 -81102 -1448 -76748
rect -2147 -81130 -1448 -81102
rect -1428 -76748 -729 -76720
rect -1428 -81102 -813 -76748
rect -749 -81102 -729 -76748
rect -1428 -81130 -729 -81102
rect -709 -76748 -10 -76720
rect -709 -81102 -94 -76748
rect -30 -81102 -10 -76748
rect -709 -81130 -10 -81102
rect 10 -76748 709 -76720
rect 10 -81102 625 -76748
rect 689 -81102 709 -76748
rect 10 -81130 709 -81102
rect 729 -76748 1428 -76720
rect 729 -81102 1344 -76748
rect 1408 -81102 1428 -76748
rect 729 -81130 1428 -81102
rect 1448 -76748 2147 -76720
rect 1448 -81102 2063 -76748
rect 2127 -81102 2147 -76748
rect 1448 -81130 2147 -81102
rect 2167 -76748 2866 -76720
rect 2167 -81102 2782 -76748
rect 2846 -81102 2866 -76748
rect 2167 -81130 2866 -81102
rect -2866 -81258 -2167 -81230
rect -2866 -85612 -2251 -81258
rect -2187 -85612 -2167 -81258
rect -2866 -85640 -2167 -85612
rect -2147 -81258 -1448 -81230
rect -2147 -85612 -1532 -81258
rect -1468 -85612 -1448 -81258
rect -2147 -85640 -1448 -85612
rect -1428 -81258 -729 -81230
rect -1428 -85612 -813 -81258
rect -749 -85612 -729 -81258
rect -1428 -85640 -729 -85612
rect -709 -81258 -10 -81230
rect -709 -85612 -94 -81258
rect -30 -85612 -10 -81258
rect -709 -85640 -10 -85612
rect 10 -81258 709 -81230
rect 10 -85612 625 -81258
rect 689 -85612 709 -81258
rect 10 -85640 709 -85612
rect 729 -81258 1428 -81230
rect 729 -85612 1344 -81258
rect 1408 -85612 1428 -81258
rect 729 -85640 1428 -85612
rect 1448 -81258 2147 -81230
rect 1448 -85612 2063 -81258
rect 2127 -85612 2147 -81258
rect 1448 -85640 2147 -85612
rect 2167 -81258 2866 -81230
rect 2167 -85612 2782 -81258
rect 2846 -85612 2866 -81258
rect 2167 -85640 2866 -85612
rect -2866 -85768 -2167 -85740
rect -2866 -90122 -2251 -85768
rect -2187 -90122 -2167 -85768
rect -2866 -90150 -2167 -90122
rect -2147 -85768 -1448 -85740
rect -2147 -90122 -1532 -85768
rect -1468 -90122 -1448 -85768
rect -2147 -90150 -1448 -90122
rect -1428 -85768 -729 -85740
rect -1428 -90122 -813 -85768
rect -749 -90122 -729 -85768
rect -1428 -90150 -729 -90122
rect -709 -85768 -10 -85740
rect -709 -90122 -94 -85768
rect -30 -90122 -10 -85768
rect -709 -90150 -10 -90122
rect 10 -85768 709 -85740
rect 10 -90122 625 -85768
rect 689 -90122 709 -85768
rect 10 -90150 709 -90122
rect 729 -85768 1428 -85740
rect 729 -90122 1344 -85768
rect 1408 -90122 1428 -85768
rect 729 -90150 1428 -90122
rect 1448 -85768 2147 -85740
rect 1448 -90122 2063 -85768
rect 2127 -90122 2147 -85768
rect 1448 -90150 2147 -90122
rect 2167 -85768 2866 -85740
rect 2167 -90122 2782 -85768
rect 2846 -90122 2866 -85768
rect 2167 -90150 2866 -90122
rect -2866 -90278 -2167 -90250
rect -2866 -94632 -2251 -90278
rect -2187 -94632 -2167 -90278
rect -2866 -94660 -2167 -94632
rect -2147 -90278 -1448 -90250
rect -2147 -94632 -1532 -90278
rect -1468 -94632 -1448 -90278
rect -2147 -94660 -1448 -94632
rect -1428 -90278 -729 -90250
rect -1428 -94632 -813 -90278
rect -749 -94632 -729 -90278
rect -1428 -94660 -729 -94632
rect -709 -90278 -10 -90250
rect -709 -94632 -94 -90278
rect -30 -94632 -10 -90278
rect -709 -94660 -10 -94632
rect 10 -90278 709 -90250
rect 10 -94632 625 -90278
rect 689 -94632 709 -90278
rect 10 -94660 709 -94632
rect 729 -90278 1428 -90250
rect 729 -94632 1344 -90278
rect 1408 -94632 1428 -90278
rect 729 -94660 1428 -94632
rect 1448 -90278 2147 -90250
rect 1448 -94632 2063 -90278
rect 2127 -94632 2147 -90278
rect 1448 -94660 2147 -94632
rect 2167 -90278 2866 -90250
rect 2167 -94632 2782 -90278
rect 2846 -94632 2866 -90278
rect 2167 -94660 2866 -94632
rect -2866 -94788 -2167 -94760
rect -2866 -99142 -2251 -94788
rect -2187 -99142 -2167 -94788
rect -2866 -99170 -2167 -99142
rect -2147 -94788 -1448 -94760
rect -2147 -99142 -1532 -94788
rect -1468 -99142 -1448 -94788
rect -2147 -99170 -1448 -99142
rect -1428 -94788 -729 -94760
rect -1428 -99142 -813 -94788
rect -749 -99142 -729 -94788
rect -1428 -99170 -729 -99142
rect -709 -94788 -10 -94760
rect -709 -99142 -94 -94788
rect -30 -99142 -10 -94788
rect -709 -99170 -10 -99142
rect 10 -94788 709 -94760
rect 10 -99142 625 -94788
rect 689 -99142 709 -94788
rect 10 -99170 709 -99142
rect 729 -94788 1428 -94760
rect 729 -99142 1344 -94788
rect 1408 -99142 1428 -94788
rect 729 -99170 1428 -99142
rect 1448 -94788 2147 -94760
rect 1448 -99142 2063 -94788
rect 2127 -99142 2147 -94788
rect 1448 -99170 2147 -99142
rect 2167 -94788 2866 -94760
rect 2167 -99142 2782 -94788
rect 2846 -99142 2866 -94788
rect 2167 -99170 2866 -99142
rect -2866 -99298 -2167 -99270
rect -2866 -103652 -2251 -99298
rect -2187 -103652 -2167 -99298
rect -2866 -103680 -2167 -103652
rect -2147 -99298 -1448 -99270
rect -2147 -103652 -1532 -99298
rect -1468 -103652 -1448 -99298
rect -2147 -103680 -1448 -103652
rect -1428 -99298 -729 -99270
rect -1428 -103652 -813 -99298
rect -749 -103652 -729 -99298
rect -1428 -103680 -729 -103652
rect -709 -99298 -10 -99270
rect -709 -103652 -94 -99298
rect -30 -103652 -10 -99298
rect -709 -103680 -10 -103652
rect 10 -99298 709 -99270
rect 10 -103652 625 -99298
rect 689 -103652 709 -99298
rect 10 -103680 709 -103652
rect 729 -99298 1428 -99270
rect 729 -103652 1344 -99298
rect 1408 -103652 1428 -99298
rect 729 -103680 1428 -103652
rect 1448 -99298 2147 -99270
rect 1448 -103652 2063 -99298
rect 2127 -103652 2147 -99298
rect 1448 -103680 2147 -103652
rect 2167 -99298 2866 -99270
rect 2167 -103652 2782 -99298
rect 2846 -103652 2866 -99298
rect 2167 -103680 2866 -103652
rect -2866 -103808 -2167 -103780
rect -2866 -108162 -2251 -103808
rect -2187 -108162 -2167 -103808
rect -2866 -108190 -2167 -108162
rect -2147 -103808 -1448 -103780
rect -2147 -108162 -1532 -103808
rect -1468 -108162 -1448 -103808
rect -2147 -108190 -1448 -108162
rect -1428 -103808 -729 -103780
rect -1428 -108162 -813 -103808
rect -749 -108162 -729 -103808
rect -1428 -108190 -729 -108162
rect -709 -103808 -10 -103780
rect -709 -108162 -94 -103808
rect -30 -108162 -10 -103808
rect -709 -108190 -10 -108162
rect 10 -103808 709 -103780
rect 10 -108162 625 -103808
rect 689 -108162 709 -103808
rect 10 -108190 709 -108162
rect 729 -103808 1428 -103780
rect 729 -108162 1344 -103808
rect 1408 -108162 1428 -103808
rect 729 -108190 1428 -108162
rect 1448 -103808 2147 -103780
rect 1448 -108162 2063 -103808
rect 2127 -108162 2147 -103808
rect 1448 -108190 2147 -108162
rect 2167 -103808 2866 -103780
rect 2167 -108162 2782 -103808
rect 2846 -108162 2866 -103808
rect 2167 -108190 2866 -108162
rect -2866 -108318 -2167 -108290
rect -2866 -112672 -2251 -108318
rect -2187 -112672 -2167 -108318
rect -2866 -112700 -2167 -112672
rect -2147 -108318 -1448 -108290
rect -2147 -112672 -1532 -108318
rect -1468 -112672 -1448 -108318
rect -2147 -112700 -1448 -112672
rect -1428 -108318 -729 -108290
rect -1428 -112672 -813 -108318
rect -749 -112672 -729 -108318
rect -1428 -112700 -729 -112672
rect -709 -108318 -10 -108290
rect -709 -112672 -94 -108318
rect -30 -112672 -10 -108318
rect -709 -112700 -10 -112672
rect 10 -108318 709 -108290
rect 10 -112672 625 -108318
rect 689 -112672 709 -108318
rect 10 -112700 709 -112672
rect 729 -108318 1428 -108290
rect 729 -112672 1344 -108318
rect 1408 -112672 1428 -108318
rect 729 -112700 1428 -112672
rect 1448 -108318 2147 -108290
rect 1448 -112672 2063 -108318
rect 2127 -112672 2147 -108318
rect 1448 -112700 2147 -112672
rect 2167 -108318 2866 -108290
rect 2167 -112672 2782 -108318
rect 2846 -112672 2866 -108318
rect 2167 -112700 2866 -112672
rect -2866 -112828 -2167 -112800
rect -2866 -117182 -2251 -112828
rect -2187 -117182 -2167 -112828
rect -2866 -117210 -2167 -117182
rect -2147 -112828 -1448 -112800
rect -2147 -117182 -1532 -112828
rect -1468 -117182 -1448 -112828
rect -2147 -117210 -1448 -117182
rect -1428 -112828 -729 -112800
rect -1428 -117182 -813 -112828
rect -749 -117182 -729 -112828
rect -1428 -117210 -729 -117182
rect -709 -112828 -10 -112800
rect -709 -117182 -94 -112828
rect -30 -117182 -10 -112828
rect -709 -117210 -10 -117182
rect 10 -112828 709 -112800
rect 10 -117182 625 -112828
rect 689 -117182 709 -112828
rect 10 -117210 709 -117182
rect 729 -112828 1428 -112800
rect 729 -117182 1344 -112828
rect 1408 -117182 1428 -112828
rect 729 -117210 1428 -117182
rect 1448 -112828 2147 -112800
rect 1448 -117182 2063 -112828
rect 2127 -117182 2147 -112828
rect 1448 -117210 2147 -117182
rect 2167 -112828 2866 -112800
rect 2167 -117182 2782 -112828
rect 2846 -117182 2866 -112828
rect 2167 -117210 2866 -117182
rect -2866 -117338 -2167 -117310
rect -2866 -121692 -2251 -117338
rect -2187 -121692 -2167 -117338
rect -2866 -121720 -2167 -121692
rect -2147 -117338 -1448 -117310
rect -2147 -121692 -1532 -117338
rect -1468 -121692 -1448 -117338
rect -2147 -121720 -1448 -121692
rect -1428 -117338 -729 -117310
rect -1428 -121692 -813 -117338
rect -749 -121692 -729 -117338
rect -1428 -121720 -729 -121692
rect -709 -117338 -10 -117310
rect -709 -121692 -94 -117338
rect -30 -121692 -10 -117338
rect -709 -121720 -10 -121692
rect 10 -117338 709 -117310
rect 10 -121692 625 -117338
rect 689 -121692 709 -117338
rect 10 -121720 709 -121692
rect 729 -117338 1428 -117310
rect 729 -121692 1344 -117338
rect 1408 -121692 1428 -117338
rect 729 -121720 1428 -121692
rect 1448 -117338 2147 -117310
rect 1448 -121692 2063 -117338
rect 2127 -121692 2147 -117338
rect 1448 -121720 2147 -121692
rect 2167 -117338 2866 -117310
rect 2167 -121692 2782 -117338
rect 2846 -121692 2866 -117338
rect 2167 -121720 2866 -121692
rect -2866 -121848 -2167 -121820
rect -2866 -126202 -2251 -121848
rect -2187 -126202 -2167 -121848
rect -2866 -126230 -2167 -126202
rect -2147 -121848 -1448 -121820
rect -2147 -126202 -1532 -121848
rect -1468 -126202 -1448 -121848
rect -2147 -126230 -1448 -126202
rect -1428 -121848 -729 -121820
rect -1428 -126202 -813 -121848
rect -749 -126202 -729 -121848
rect -1428 -126230 -729 -126202
rect -709 -121848 -10 -121820
rect -709 -126202 -94 -121848
rect -30 -126202 -10 -121848
rect -709 -126230 -10 -126202
rect 10 -121848 709 -121820
rect 10 -126202 625 -121848
rect 689 -126202 709 -121848
rect 10 -126230 709 -126202
rect 729 -121848 1428 -121820
rect 729 -126202 1344 -121848
rect 1408 -126202 1428 -121848
rect 729 -126230 1428 -126202
rect 1448 -121848 2147 -121820
rect 1448 -126202 2063 -121848
rect 2127 -126202 2147 -121848
rect 1448 -126230 2147 -126202
rect 2167 -121848 2866 -121820
rect 2167 -126202 2782 -121848
rect 2846 -126202 2866 -121848
rect 2167 -126230 2866 -126202
rect -2866 -126358 -2167 -126330
rect -2866 -130712 -2251 -126358
rect -2187 -130712 -2167 -126358
rect -2866 -130740 -2167 -130712
rect -2147 -126358 -1448 -126330
rect -2147 -130712 -1532 -126358
rect -1468 -130712 -1448 -126358
rect -2147 -130740 -1448 -130712
rect -1428 -126358 -729 -126330
rect -1428 -130712 -813 -126358
rect -749 -130712 -729 -126358
rect -1428 -130740 -729 -130712
rect -709 -126358 -10 -126330
rect -709 -130712 -94 -126358
rect -30 -130712 -10 -126358
rect -709 -130740 -10 -130712
rect 10 -126358 709 -126330
rect 10 -130712 625 -126358
rect 689 -130712 709 -126358
rect 10 -130740 709 -130712
rect 729 -126358 1428 -126330
rect 729 -130712 1344 -126358
rect 1408 -130712 1428 -126358
rect 729 -130740 1428 -130712
rect 1448 -126358 2147 -126330
rect 1448 -130712 2063 -126358
rect 2127 -130712 2147 -126358
rect 1448 -130740 2147 -130712
rect 2167 -126358 2866 -126330
rect 2167 -130712 2782 -126358
rect 2846 -130712 2866 -126358
rect 2167 -130740 2866 -130712
rect -2866 -130868 -2167 -130840
rect -2866 -135222 -2251 -130868
rect -2187 -135222 -2167 -130868
rect -2866 -135250 -2167 -135222
rect -2147 -130868 -1448 -130840
rect -2147 -135222 -1532 -130868
rect -1468 -135222 -1448 -130868
rect -2147 -135250 -1448 -135222
rect -1428 -130868 -729 -130840
rect -1428 -135222 -813 -130868
rect -749 -135222 -729 -130868
rect -1428 -135250 -729 -135222
rect -709 -130868 -10 -130840
rect -709 -135222 -94 -130868
rect -30 -135222 -10 -130868
rect -709 -135250 -10 -135222
rect 10 -130868 709 -130840
rect 10 -135222 625 -130868
rect 689 -135222 709 -130868
rect 10 -135250 709 -135222
rect 729 -130868 1428 -130840
rect 729 -135222 1344 -130868
rect 1408 -135222 1428 -130868
rect 729 -135250 1428 -135222
rect 1448 -130868 2147 -130840
rect 1448 -135222 2063 -130868
rect 2127 -135222 2147 -130868
rect 1448 -135250 2147 -135222
rect 2167 -130868 2866 -130840
rect 2167 -135222 2782 -130868
rect 2846 -135222 2866 -130868
rect 2167 -135250 2866 -135222
rect -2866 -135378 -2167 -135350
rect -2866 -139732 -2251 -135378
rect -2187 -139732 -2167 -135378
rect -2866 -139760 -2167 -139732
rect -2147 -135378 -1448 -135350
rect -2147 -139732 -1532 -135378
rect -1468 -139732 -1448 -135378
rect -2147 -139760 -1448 -139732
rect -1428 -135378 -729 -135350
rect -1428 -139732 -813 -135378
rect -749 -139732 -729 -135378
rect -1428 -139760 -729 -139732
rect -709 -135378 -10 -135350
rect -709 -139732 -94 -135378
rect -30 -139732 -10 -135378
rect -709 -139760 -10 -139732
rect 10 -135378 709 -135350
rect 10 -139732 625 -135378
rect 689 -139732 709 -135378
rect 10 -139760 709 -139732
rect 729 -135378 1428 -135350
rect 729 -139732 1344 -135378
rect 1408 -139732 1428 -135378
rect 729 -139760 1428 -139732
rect 1448 -135378 2147 -135350
rect 1448 -139732 2063 -135378
rect 2127 -139732 2147 -135378
rect 1448 -139760 2147 -139732
rect 2167 -135378 2866 -135350
rect 2167 -139732 2782 -135378
rect 2846 -139732 2866 -135378
rect 2167 -139760 2866 -139732
rect -2866 -139888 -2167 -139860
rect -2866 -144242 -2251 -139888
rect -2187 -144242 -2167 -139888
rect -2866 -144270 -2167 -144242
rect -2147 -139888 -1448 -139860
rect -2147 -144242 -1532 -139888
rect -1468 -144242 -1448 -139888
rect -2147 -144270 -1448 -144242
rect -1428 -139888 -729 -139860
rect -1428 -144242 -813 -139888
rect -749 -144242 -729 -139888
rect -1428 -144270 -729 -144242
rect -709 -139888 -10 -139860
rect -709 -144242 -94 -139888
rect -30 -144242 -10 -139888
rect -709 -144270 -10 -144242
rect 10 -139888 709 -139860
rect 10 -144242 625 -139888
rect 689 -144242 709 -139888
rect 10 -144270 709 -144242
rect 729 -139888 1428 -139860
rect 729 -144242 1344 -139888
rect 1408 -144242 1428 -139888
rect 729 -144270 1428 -144242
rect 1448 -139888 2147 -139860
rect 1448 -144242 2063 -139888
rect 2127 -144242 2147 -139888
rect 1448 -144270 2147 -144242
rect 2167 -139888 2866 -139860
rect 2167 -144242 2782 -139888
rect 2846 -144242 2866 -139888
rect 2167 -144270 2866 -144242
<< via3 >>
rect -2251 139888 -2187 144242
rect -1532 139888 -1468 144242
rect -813 139888 -749 144242
rect -94 139888 -30 144242
rect 625 139888 689 144242
rect 1344 139888 1408 144242
rect 2063 139888 2127 144242
rect 2782 139888 2846 144242
rect -2251 135378 -2187 139732
rect -1532 135378 -1468 139732
rect -813 135378 -749 139732
rect -94 135378 -30 139732
rect 625 135378 689 139732
rect 1344 135378 1408 139732
rect 2063 135378 2127 139732
rect 2782 135378 2846 139732
rect -2251 130868 -2187 135222
rect -1532 130868 -1468 135222
rect -813 130868 -749 135222
rect -94 130868 -30 135222
rect 625 130868 689 135222
rect 1344 130868 1408 135222
rect 2063 130868 2127 135222
rect 2782 130868 2846 135222
rect -2251 126358 -2187 130712
rect -1532 126358 -1468 130712
rect -813 126358 -749 130712
rect -94 126358 -30 130712
rect 625 126358 689 130712
rect 1344 126358 1408 130712
rect 2063 126358 2127 130712
rect 2782 126358 2846 130712
rect -2251 121848 -2187 126202
rect -1532 121848 -1468 126202
rect -813 121848 -749 126202
rect -94 121848 -30 126202
rect 625 121848 689 126202
rect 1344 121848 1408 126202
rect 2063 121848 2127 126202
rect 2782 121848 2846 126202
rect -2251 117338 -2187 121692
rect -1532 117338 -1468 121692
rect -813 117338 -749 121692
rect -94 117338 -30 121692
rect 625 117338 689 121692
rect 1344 117338 1408 121692
rect 2063 117338 2127 121692
rect 2782 117338 2846 121692
rect -2251 112828 -2187 117182
rect -1532 112828 -1468 117182
rect -813 112828 -749 117182
rect -94 112828 -30 117182
rect 625 112828 689 117182
rect 1344 112828 1408 117182
rect 2063 112828 2127 117182
rect 2782 112828 2846 117182
rect -2251 108318 -2187 112672
rect -1532 108318 -1468 112672
rect -813 108318 -749 112672
rect -94 108318 -30 112672
rect 625 108318 689 112672
rect 1344 108318 1408 112672
rect 2063 108318 2127 112672
rect 2782 108318 2846 112672
rect -2251 103808 -2187 108162
rect -1532 103808 -1468 108162
rect -813 103808 -749 108162
rect -94 103808 -30 108162
rect 625 103808 689 108162
rect 1344 103808 1408 108162
rect 2063 103808 2127 108162
rect 2782 103808 2846 108162
rect -2251 99298 -2187 103652
rect -1532 99298 -1468 103652
rect -813 99298 -749 103652
rect -94 99298 -30 103652
rect 625 99298 689 103652
rect 1344 99298 1408 103652
rect 2063 99298 2127 103652
rect 2782 99298 2846 103652
rect -2251 94788 -2187 99142
rect -1532 94788 -1468 99142
rect -813 94788 -749 99142
rect -94 94788 -30 99142
rect 625 94788 689 99142
rect 1344 94788 1408 99142
rect 2063 94788 2127 99142
rect 2782 94788 2846 99142
rect -2251 90278 -2187 94632
rect -1532 90278 -1468 94632
rect -813 90278 -749 94632
rect -94 90278 -30 94632
rect 625 90278 689 94632
rect 1344 90278 1408 94632
rect 2063 90278 2127 94632
rect 2782 90278 2846 94632
rect -2251 85768 -2187 90122
rect -1532 85768 -1468 90122
rect -813 85768 -749 90122
rect -94 85768 -30 90122
rect 625 85768 689 90122
rect 1344 85768 1408 90122
rect 2063 85768 2127 90122
rect 2782 85768 2846 90122
rect -2251 81258 -2187 85612
rect -1532 81258 -1468 85612
rect -813 81258 -749 85612
rect -94 81258 -30 85612
rect 625 81258 689 85612
rect 1344 81258 1408 85612
rect 2063 81258 2127 85612
rect 2782 81258 2846 85612
rect -2251 76748 -2187 81102
rect -1532 76748 -1468 81102
rect -813 76748 -749 81102
rect -94 76748 -30 81102
rect 625 76748 689 81102
rect 1344 76748 1408 81102
rect 2063 76748 2127 81102
rect 2782 76748 2846 81102
rect -2251 72238 -2187 76592
rect -1532 72238 -1468 76592
rect -813 72238 -749 76592
rect -94 72238 -30 76592
rect 625 72238 689 76592
rect 1344 72238 1408 76592
rect 2063 72238 2127 76592
rect 2782 72238 2846 76592
rect -2251 67728 -2187 72082
rect -1532 67728 -1468 72082
rect -813 67728 -749 72082
rect -94 67728 -30 72082
rect 625 67728 689 72082
rect 1344 67728 1408 72082
rect 2063 67728 2127 72082
rect 2782 67728 2846 72082
rect -2251 63218 -2187 67572
rect -1532 63218 -1468 67572
rect -813 63218 -749 67572
rect -94 63218 -30 67572
rect 625 63218 689 67572
rect 1344 63218 1408 67572
rect 2063 63218 2127 67572
rect 2782 63218 2846 67572
rect -2251 58708 -2187 63062
rect -1532 58708 -1468 63062
rect -813 58708 -749 63062
rect -94 58708 -30 63062
rect 625 58708 689 63062
rect 1344 58708 1408 63062
rect 2063 58708 2127 63062
rect 2782 58708 2846 63062
rect -2251 54198 -2187 58552
rect -1532 54198 -1468 58552
rect -813 54198 -749 58552
rect -94 54198 -30 58552
rect 625 54198 689 58552
rect 1344 54198 1408 58552
rect 2063 54198 2127 58552
rect 2782 54198 2846 58552
rect -2251 49688 -2187 54042
rect -1532 49688 -1468 54042
rect -813 49688 -749 54042
rect -94 49688 -30 54042
rect 625 49688 689 54042
rect 1344 49688 1408 54042
rect 2063 49688 2127 54042
rect 2782 49688 2846 54042
rect -2251 45178 -2187 49532
rect -1532 45178 -1468 49532
rect -813 45178 -749 49532
rect -94 45178 -30 49532
rect 625 45178 689 49532
rect 1344 45178 1408 49532
rect 2063 45178 2127 49532
rect 2782 45178 2846 49532
rect -2251 40668 -2187 45022
rect -1532 40668 -1468 45022
rect -813 40668 -749 45022
rect -94 40668 -30 45022
rect 625 40668 689 45022
rect 1344 40668 1408 45022
rect 2063 40668 2127 45022
rect 2782 40668 2846 45022
rect -2251 36158 -2187 40512
rect -1532 36158 -1468 40512
rect -813 36158 -749 40512
rect -94 36158 -30 40512
rect 625 36158 689 40512
rect 1344 36158 1408 40512
rect 2063 36158 2127 40512
rect 2782 36158 2846 40512
rect -2251 31648 -2187 36002
rect -1532 31648 -1468 36002
rect -813 31648 -749 36002
rect -94 31648 -30 36002
rect 625 31648 689 36002
rect 1344 31648 1408 36002
rect 2063 31648 2127 36002
rect 2782 31648 2846 36002
rect -2251 27138 -2187 31492
rect -1532 27138 -1468 31492
rect -813 27138 -749 31492
rect -94 27138 -30 31492
rect 625 27138 689 31492
rect 1344 27138 1408 31492
rect 2063 27138 2127 31492
rect 2782 27138 2846 31492
rect -2251 22628 -2187 26982
rect -1532 22628 -1468 26982
rect -813 22628 -749 26982
rect -94 22628 -30 26982
rect 625 22628 689 26982
rect 1344 22628 1408 26982
rect 2063 22628 2127 26982
rect 2782 22628 2846 26982
rect -2251 18118 -2187 22472
rect -1532 18118 -1468 22472
rect -813 18118 -749 22472
rect -94 18118 -30 22472
rect 625 18118 689 22472
rect 1344 18118 1408 22472
rect 2063 18118 2127 22472
rect 2782 18118 2846 22472
rect -2251 13608 -2187 17962
rect -1532 13608 -1468 17962
rect -813 13608 -749 17962
rect -94 13608 -30 17962
rect 625 13608 689 17962
rect 1344 13608 1408 17962
rect 2063 13608 2127 17962
rect 2782 13608 2846 17962
rect -2251 9098 -2187 13452
rect -1532 9098 -1468 13452
rect -813 9098 -749 13452
rect -94 9098 -30 13452
rect 625 9098 689 13452
rect 1344 9098 1408 13452
rect 2063 9098 2127 13452
rect 2782 9098 2846 13452
rect -2251 4588 -2187 8942
rect -1532 4588 -1468 8942
rect -813 4588 -749 8942
rect -94 4588 -30 8942
rect 625 4588 689 8942
rect 1344 4588 1408 8942
rect 2063 4588 2127 8942
rect 2782 4588 2846 8942
rect -2251 78 -2187 4432
rect -1532 78 -1468 4432
rect -813 78 -749 4432
rect -94 78 -30 4432
rect 625 78 689 4432
rect 1344 78 1408 4432
rect 2063 78 2127 4432
rect 2782 78 2846 4432
rect -2251 -4432 -2187 -78
rect -1532 -4432 -1468 -78
rect -813 -4432 -749 -78
rect -94 -4432 -30 -78
rect 625 -4432 689 -78
rect 1344 -4432 1408 -78
rect 2063 -4432 2127 -78
rect 2782 -4432 2846 -78
rect -2251 -8942 -2187 -4588
rect -1532 -8942 -1468 -4588
rect -813 -8942 -749 -4588
rect -94 -8942 -30 -4588
rect 625 -8942 689 -4588
rect 1344 -8942 1408 -4588
rect 2063 -8942 2127 -4588
rect 2782 -8942 2846 -4588
rect -2251 -13452 -2187 -9098
rect -1532 -13452 -1468 -9098
rect -813 -13452 -749 -9098
rect -94 -13452 -30 -9098
rect 625 -13452 689 -9098
rect 1344 -13452 1408 -9098
rect 2063 -13452 2127 -9098
rect 2782 -13452 2846 -9098
rect -2251 -17962 -2187 -13608
rect -1532 -17962 -1468 -13608
rect -813 -17962 -749 -13608
rect -94 -17962 -30 -13608
rect 625 -17962 689 -13608
rect 1344 -17962 1408 -13608
rect 2063 -17962 2127 -13608
rect 2782 -17962 2846 -13608
rect -2251 -22472 -2187 -18118
rect -1532 -22472 -1468 -18118
rect -813 -22472 -749 -18118
rect -94 -22472 -30 -18118
rect 625 -22472 689 -18118
rect 1344 -22472 1408 -18118
rect 2063 -22472 2127 -18118
rect 2782 -22472 2846 -18118
rect -2251 -26982 -2187 -22628
rect -1532 -26982 -1468 -22628
rect -813 -26982 -749 -22628
rect -94 -26982 -30 -22628
rect 625 -26982 689 -22628
rect 1344 -26982 1408 -22628
rect 2063 -26982 2127 -22628
rect 2782 -26982 2846 -22628
rect -2251 -31492 -2187 -27138
rect -1532 -31492 -1468 -27138
rect -813 -31492 -749 -27138
rect -94 -31492 -30 -27138
rect 625 -31492 689 -27138
rect 1344 -31492 1408 -27138
rect 2063 -31492 2127 -27138
rect 2782 -31492 2846 -27138
rect -2251 -36002 -2187 -31648
rect -1532 -36002 -1468 -31648
rect -813 -36002 -749 -31648
rect -94 -36002 -30 -31648
rect 625 -36002 689 -31648
rect 1344 -36002 1408 -31648
rect 2063 -36002 2127 -31648
rect 2782 -36002 2846 -31648
rect -2251 -40512 -2187 -36158
rect -1532 -40512 -1468 -36158
rect -813 -40512 -749 -36158
rect -94 -40512 -30 -36158
rect 625 -40512 689 -36158
rect 1344 -40512 1408 -36158
rect 2063 -40512 2127 -36158
rect 2782 -40512 2846 -36158
rect -2251 -45022 -2187 -40668
rect -1532 -45022 -1468 -40668
rect -813 -45022 -749 -40668
rect -94 -45022 -30 -40668
rect 625 -45022 689 -40668
rect 1344 -45022 1408 -40668
rect 2063 -45022 2127 -40668
rect 2782 -45022 2846 -40668
rect -2251 -49532 -2187 -45178
rect -1532 -49532 -1468 -45178
rect -813 -49532 -749 -45178
rect -94 -49532 -30 -45178
rect 625 -49532 689 -45178
rect 1344 -49532 1408 -45178
rect 2063 -49532 2127 -45178
rect 2782 -49532 2846 -45178
rect -2251 -54042 -2187 -49688
rect -1532 -54042 -1468 -49688
rect -813 -54042 -749 -49688
rect -94 -54042 -30 -49688
rect 625 -54042 689 -49688
rect 1344 -54042 1408 -49688
rect 2063 -54042 2127 -49688
rect 2782 -54042 2846 -49688
rect -2251 -58552 -2187 -54198
rect -1532 -58552 -1468 -54198
rect -813 -58552 -749 -54198
rect -94 -58552 -30 -54198
rect 625 -58552 689 -54198
rect 1344 -58552 1408 -54198
rect 2063 -58552 2127 -54198
rect 2782 -58552 2846 -54198
rect -2251 -63062 -2187 -58708
rect -1532 -63062 -1468 -58708
rect -813 -63062 -749 -58708
rect -94 -63062 -30 -58708
rect 625 -63062 689 -58708
rect 1344 -63062 1408 -58708
rect 2063 -63062 2127 -58708
rect 2782 -63062 2846 -58708
rect -2251 -67572 -2187 -63218
rect -1532 -67572 -1468 -63218
rect -813 -67572 -749 -63218
rect -94 -67572 -30 -63218
rect 625 -67572 689 -63218
rect 1344 -67572 1408 -63218
rect 2063 -67572 2127 -63218
rect 2782 -67572 2846 -63218
rect -2251 -72082 -2187 -67728
rect -1532 -72082 -1468 -67728
rect -813 -72082 -749 -67728
rect -94 -72082 -30 -67728
rect 625 -72082 689 -67728
rect 1344 -72082 1408 -67728
rect 2063 -72082 2127 -67728
rect 2782 -72082 2846 -67728
rect -2251 -76592 -2187 -72238
rect -1532 -76592 -1468 -72238
rect -813 -76592 -749 -72238
rect -94 -76592 -30 -72238
rect 625 -76592 689 -72238
rect 1344 -76592 1408 -72238
rect 2063 -76592 2127 -72238
rect 2782 -76592 2846 -72238
rect -2251 -81102 -2187 -76748
rect -1532 -81102 -1468 -76748
rect -813 -81102 -749 -76748
rect -94 -81102 -30 -76748
rect 625 -81102 689 -76748
rect 1344 -81102 1408 -76748
rect 2063 -81102 2127 -76748
rect 2782 -81102 2846 -76748
rect -2251 -85612 -2187 -81258
rect -1532 -85612 -1468 -81258
rect -813 -85612 -749 -81258
rect -94 -85612 -30 -81258
rect 625 -85612 689 -81258
rect 1344 -85612 1408 -81258
rect 2063 -85612 2127 -81258
rect 2782 -85612 2846 -81258
rect -2251 -90122 -2187 -85768
rect -1532 -90122 -1468 -85768
rect -813 -90122 -749 -85768
rect -94 -90122 -30 -85768
rect 625 -90122 689 -85768
rect 1344 -90122 1408 -85768
rect 2063 -90122 2127 -85768
rect 2782 -90122 2846 -85768
rect -2251 -94632 -2187 -90278
rect -1532 -94632 -1468 -90278
rect -813 -94632 -749 -90278
rect -94 -94632 -30 -90278
rect 625 -94632 689 -90278
rect 1344 -94632 1408 -90278
rect 2063 -94632 2127 -90278
rect 2782 -94632 2846 -90278
rect -2251 -99142 -2187 -94788
rect -1532 -99142 -1468 -94788
rect -813 -99142 -749 -94788
rect -94 -99142 -30 -94788
rect 625 -99142 689 -94788
rect 1344 -99142 1408 -94788
rect 2063 -99142 2127 -94788
rect 2782 -99142 2846 -94788
rect -2251 -103652 -2187 -99298
rect -1532 -103652 -1468 -99298
rect -813 -103652 -749 -99298
rect -94 -103652 -30 -99298
rect 625 -103652 689 -99298
rect 1344 -103652 1408 -99298
rect 2063 -103652 2127 -99298
rect 2782 -103652 2846 -99298
rect -2251 -108162 -2187 -103808
rect -1532 -108162 -1468 -103808
rect -813 -108162 -749 -103808
rect -94 -108162 -30 -103808
rect 625 -108162 689 -103808
rect 1344 -108162 1408 -103808
rect 2063 -108162 2127 -103808
rect 2782 -108162 2846 -103808
rect -2251 -112672 -2187 -108318
rect -1532 -112672 -1468 -108318
rect -813 -112672 -749 -108318
rect -94 -112672 -30 -108318
rect 625 -112672 689 -108318
rect 1344 -112672 1408 -108318
rect 2063 -112672 2127 -108318
rect 2782 -112672 2846 -108318
rect -2251 -117182 -2187 -112828
rect -1532 -117182 -1468 -112828
rect -813 -117182 -749 -112828
rect -94 -117182 -30 -112828
rect 625 -117182 689 -112828
rect 1344 -117182 1408 -112828
rect 2063 -117182 2127 -112828
rect 2782 -117182 2846 -112828
rect -2251 -121692 -2187 -117338
rect -1532 -121692 -1468 -117338
rect -813 -121692 -749 -117338
rect -94 -121692 -30 -117338
rect 625 -121692 689 -117338
rect 1344 -121692 1408 -117338
rect 2063 -121692 2127 -117338
rect 2782 -121692 2846 -117338
rect -2251 -126202 -2187 -121848
rect -1532 -126202 -1468 -121848
rect -813 -126202 -749 -121848
rect -94 -126202 -30 -121848
rect 625 -126202 689 -121848
rect 1344 -126202 1408 -121848
rect 2063 -126202 2127 -121848
rect 2782 -126202 2846 -121848
rect -2251 -130712 -2187 -126358
rect -1532 -130712 -1468 -126358
rect -813 -130712 -749 -126358
rect -94 -130712 -30 -126358
rect 625 -130712 689 -126358
rect 1344 -130712 1408 -126358
rect 2063 -130712 2127 -126358
rect 2782 -130712 2846 -126358
rect -2251 -135222 -2187 -130868
rect -1532 -135222 -1468 -130868
rect -813 -135222 -749 -130868
rect -94 -135222 -30 -130868
rect 625 -135222 689 -130868
rect 1344 -135222 1408 -130868
rect 2063 -135222 2127 -130868
rect 2782 -135222 2846 -130868
rect -2251 -139732 -2187 -135378
rect -1532 -139732 -1468 -135378
rect -813 -139732 -749 -135378
rect -94 -139732 -30 -135378
rect 625 -139732 689 -135378
rect 1344 -139732 1408 -135378
rect 2063 -139732 2127 -135378
rect 2782 -139732 2846 -135378
rect -2251 -144242 -2187 -139888
rect -1532 -144242 -1468 -139888
rect -813 -144242 -749 -139888
rect -94 -144242 -30 -139888
rect 625 -144242 689 -139888
rect 1344 -144242 1408 -139888
rect 2063 -144242 2127 -139888
rect 2782 -144242 2846 -139888
<< mimcap >>
rect -2766 144130 -2366 144170
rect -2766 140000 -2726 144130
rect -2406 140000 -2366 144130
rect -2766 139960 -2366 140000
rect -2047 144130 -1647 144170
rect -2047 140000 -2007 144130
rect -1687 140000 -1647 144130
rect -2047 139960 -1647 140000
rect -1328 144130 -928 144170
rect -1328 140000 -1288 144130
rect -968 140000 -928 144130
rect -1328 139960 -928 140000
rect -609 144130 -209 144170
rect -609 140000 -569 144130
rect -249 140000 -209 144130
rect -609 139960 -209 140000
rect 110 144130 510 144170
rect 110 140000 150 144130
rect 470 140000 510 144130
rect 110 139960 510 140000
rect 829 144130 1229 144170
rect 829 140000 869 144130
rect 1189 140000 1229 144130
rect 829 139960 1229 140000
rect 1548 144130 1948 144170
rect 1548 140000 1588 144130
rect 1908 140000 1948 144130
rect 1548 139960 1948 140000
rect 2267 144130 2667 144170
rect 2267 140000 2307 144130
rect 2627 140000 2667 144130
rect 2267 139960 2667 140000
rect -2766 139620 -2366 139660
rect -2766 135490 -2726 139620
rect -2406 135490 -2366 139620
rect -2766 135450 -2366 135490
rect -2047 139620 -1647 139660
rect -2047 135490 -2007 139620
rect -1687 135490 -1647 139620
rect -2047 135450 -1647 135490
rect -1328 139620 -928 139660
rect -1328 135490 -1288 139620
rect -968 135490 -928 139620
rect -1328 135450 -928 135490
rect -609 139620 -209 139660
rect -609 135490 -569 139620
rect -249 135490 -209 139620
rect -609 135450 -209 135490
rect 110 139620 510 139660
rect 110 135490 150 139620
rect 470 135490 510 139620
rect 110 135450 510 135490
rect 829 139620 1229 139660
rect 829 135490 869 139620
rect 1189 135490 1229 139620
rect 829 135450 1229 135490
rect 1548 139620 1948 139660
rect 1548 135490 1588 139620
rect 1908 135490 1948 139620
rect 1548 135450 1948 135490
rect 2267 139620 2667 139660
rect 2267 135490 2307 139620
rect 2627 135490 2667 139620
rect 2267 135450 2667 135490
rect -2766 135110 -2366 135150
rect -2766 130980 -2726 135110
rect -2406 130980 -2366 135110
rect -2766 130940 -2366 130980
rect -2047 135110 -1647 135150
rect -2047 130980 -2007 135110
rect -1687 130980 -1647 135110
rect -2047 130940 -1647 130980
rect -1328 135110 -928 135150
rect -1328 130980 -1288 135110
rect -968 130980 -928 135110
rect -1328 130940 -928 130980
rect -609 135110 -209 135150
rect -609 130980 -569 135110
rect -249 130980 -209 135110
rect -609 130940 -209 130980
rect 110 135110 510 135150
rect 110 130980 150 135110
rect 470 130980 510 135110
rect 110 130940 510 130980
rect 829 135110 1229 135150
rect 829 130980 869 135110
rect 1189 130980 1229 135110
rect 829 130940 1229 130980
rect 1548 135110 1948 135150
rect 1548 130980 1588 135110
rect 1908 130980 1948 135110
rect 1548 130940 1948 130980
rect 2267 135110 2667 135150
rect 2267 130980 2307 135110
rect 2627 130980 2667 135110
rect 2267 130940 2667 130980
rect -2766 130600 -2366 130640
rect -2766 126470 -2726 130600
rect -2406 126470 -2366 130600
rect -2766 126430 -2366 126470
rect -2047 130600 -1647 130640
rect -2047 126470 -2007 130600
rect -1687 126470 -1647 130600
rect -2047 126430 -1647 126470
rect -1328 130600 -928 130640
rect -1328 126470 -1288 130600
rect -968 126470 -928 130600
rect -1328 126430 -928 126470
rect -609 130600 -209 130640
rect -609 126470 -569 130600
rect -249 126470 -209 130600
rect -609 126430 -209 126470
rect 110 130600 510 130640
rect 110 126470 150 130600
rect 470 126470 510 130600
rect 110 126430 510 126470
rect 829 130600 1229 130640
rect 829 126470 869 130600
rect 1189 126470 1229 130600
rect 829 126430 1229 126470
rect 1548 130600 1948 130640
rect 1548 126470 1588 130600
rect 1908 126470 1948 130600
rect 1548 126430 1948 126470
rect 2267 130600 2667 130640
rect 2267 126470 2307 130600
rect 2627 126470 2667 130600
rect 2267 126430 2667 126470
rect -2766 126090 -2366 126130
rect -2766 121960 -2726 126090
rect -2406 121960 -2366 126090
rect -2766 121920 -2366 121960
rect -2047 126090 -1647 126130
rect -2047 121960 -2007 126090
rect -1687 121960 -1647 126090
rect -2047 121920 -1647 121960
rect -1328 126090 -928 126130
rect -1328 121960 -1288 126090
rect -968 121960 -928 126090
rect -1328 121920 -928 121960
rect -609 126090 -209 126130
rect -609 121960 -569 126090
rect -249 121960 -209 126090
rect -609 121920 -209 121960
rect 110 126090 510 126130
rect 110 121960 150 126090
rect 470 121960 510 126090
rect 110 121920 510 121960
rect 829 126090 1229 126130
rect 829 121960 869 126090
rect 1189 121960 1229 126090
rect 829 121920 1229 121960
rect 1548 126090 1948 126130
rect 1548 121960 1588 126090
rect 1908 121960 1948 126090
rect 1548 121920 1948 121960
rect 2267 126090 2667 126130
rect 2267 121960 2307 126090
rect 2627 121960 2667 126090
rect 2267 121920 2667 121960
rect -2766 121580 -2366 121620
rect -2766 117450 -2726 121580
rect -2406 117450 -2366 121580
rect -2766 117410 -2366 117450
rect -2047 121580 -1647 121620
rect -2047 117450 -2007 121580
rect -1687 117450 -1647 121580
rect -2047 117410 -1647 117450
rect -1328 121580 -928 121620
rect -1328 117450 -1288 121580
rect -968 117450 -928 121580
rect -1328 117410 -928 117450
rect -609 121580 -209 121620
rect -609 117450 -569 121580
rect -249 117450 -209 121580
rect -609 117410 -209 117450
rect 110 121580 510 121620
rect 110 117450 150 121580
rect 470 117450 510 121580
rect 110 117410 510 117450
rect 829 121580 1229 121620
rect 829 117450 869 121580
rect 1189 117450 1229 121580
rect 829 117410 1229 117450
rect 1548 121580 1948 121620
rect 1548 117450 1588 121580
rect 1908 117450 1948 121580
rect 1548 117410 1948 117450
rect 2267 121580 2667 121620
rect 2267 117450 2307 121580
rect 2627 117450 2667 121580
rect 2267 117410 2667 117450
rect -2766 117070 -2366 117110
rect -2766 112940 -2726 117070
rect -2406 112940 -2366 117070
rect -2766 112900 -2366 112940
rect -2047 117070 -1647 117110
rect -2047 112940 -2007 117070
rect -1687 112940 -1647 117070
rect -2047 112900 -1647 112940
rect -1328 117070 -928 117110
rect -1328 112940 -1288 117070
rect -968 112940 -928 117070
rect -1328 112900 -928 112940
rect -609 117070 -209 117110
rect -609 112940 -569 117070
rect -249 112940 -209 117070
rect -609 112900 -209 112940
rect 110 117070 510 117110
rect 110 112940 150 117070
rect 470 112940 510 117070
rect 110 112900 510 112940
rect 829 117070 1229 117110
rect 829 112940 869 117070
rect 1189 112940 1229 117070
rect 829 112900 1229 112940
rect 1548 117070 1948 117110
rect 1548 112940 1588 117070
rect 1908 112940 1948 117070
rect 1548 112900 1948 112940
rect 2267 117070 2667 117110
rect 2267 112940 2307 117070
rect 2627 112940 2667 117070
rect 2267 112900 2667 112940
rect -2766 112560 -2366 112600
rect -2766 108430 -2726 112560
rect -2406 108430 -2366 112560
rect -2766 108390 -2366 108430
rect -2047 112560 -1647 112600
rect -2047 108430 -2007 112560
rect -1687 108430 -1647 112560
rect -2047 108390 -1647 108430
rect -1328 112560 -928 112600
rect -1328 108430 -1288 112560
rect -968 108430 -928 112560
rect -1328 108390 -928 108430
rect -609 112560 -209 112600
rect -609 108430 -569 112560
rect -249 108430 -209 112560
rect -609 108390 -209 108430
rect 110 112560 510 112600
rect 110 108430 150 112560
rect 470 108430 510 112560
rect 110 108390 510 108430
rect 829 112560 1229 112600
rect 829 108430 869 112560
rect 1189 108430 1229 112560
rect 829 108390 1229 108430
rect 1548 112560 1948 112600
rect 1548 108430 1588 112560
rect 1908 108430 1948 112560
rect 1548 108390 1948 108430
rect 2267 112560 2667 112600
rect 2267 108430 2307 112560
rect 2627 108430 2667 112560
rect 2267 108390 2667 108430
rect -2766 108050 -2366 108090
rect -2766 103920 -2726 108050
rect -2406 103920 -2366 108050
rect -2766 103880 -2366 103920
rect -2047 108050 -1647 108090
rect -2047 103920 -2007 108050
rect -1687 103920 -1647 108050
rect -2047 103880 -1647 103920
rect -1328 108050 -928 108090
rect -1328 103920 -1288 108050
rect -968 103920 -928 108050
rect -1328 103880 -928 103920
rect -609 108050 -209 108090
rect -609 103920 -569 108050
rect -249 103920 -209 108050
rect -609 103880 -209 103920
rect 110 108050 510 108090
rect 110 103920 150 108050
rect 470 103920 510 108050
rect 110 103880 510 103920
rect 829 108050 1229 108090
rect 829 103920 869 108050
rect 1189 103920 1229 108050
rect 829 103880 1229 103920
rect 1548 108050 1948 108090
rect 1548 103920 1588 108050
rect 1908 103920 1948 108050
rect 1548 103880 1948 103920
rect 2267 108050 2667 108090
rect 2267 103920 2307 108050
rect 2627 103920 2667 108050
rect 2267 103880 2667 103920
rect -2766 103540 -2366 103580
rect -2766 99410 -2726 103540
rect -2406 99410 -2366 103540
rect -2766 99370 -2366 99410
rect -2047 103540 -1647 103580
rect -2047 99410 -2007 103540
rect -1687 99410 -1647 103540
rect -2047 99370 -1647 99410
rect -1328 103540 -928 103580
rect -1328 99410 -1288 103540
rect -968 99410 -928 103540
rect -1328 99370 -928 99410
rect -609 103540 -209 103580
rect -609 99410 -569 103540
rect -249 99410 -209 103540
rect -609 99370 -209 99410
rect 110 103540 510 103580
rect 110 99410 150 103540
rect 470 99410 510 103540
rect 110 99370 510 99410
rect 829 103540 1229 103580
rect 829 99410 869 103540
rect 1189 99410 1229 103540
rect 829 99370 1229 99410
rect 1548 103540 1948 103580
rect 1548 99410 1588 103540
rect 1908 99410 1948 103540
rect 1548 99370 1948 99410
rect 2267 103540 2667 103580
rect 2267 99410 2307 103540
rect 2627 99410 2667 103540
rect 2267 99370 2667 99410
rect -2766 99030 -2366 99070
rect -2766 94900 -2726 99030
rect -2406 94900 -2366 99030
rect -2766 94860 -2366 94900
rect -2047 99030 -1647 99070
rect -2047 94900 -2007 99030
rect -1687 94900 -1647 99030
rect -2047 94860 -1647 94900
rect -1328 99030 -928 99070
rect -1328 94900 -1288 99030
rect -968 94900 -928 99030
rect -1328 94860 -928 94900
rect -609 99030 -209 99070
rect -609 94900 -569 99030
rect -249 94900 -209 99030
rect -609 94860 -209 94900
rect 110 99030 510 99070
rect 110 94900 150 99030
rect 470 94900 510 99030
rect 110 94860 510 94900
rect 829 99030 1229 99070
rect 829 94900 869 99030
rect 1189 94900 1229 99030
rect 829 94860 1229 94900
rect 1548 99030 1948 99070
rect 1548 94900 1588 99030
rect 1908 94900 1948 99030
rect 1548 94860 1948 94900
rect 2267 99030 2667 99070
rect 2267 94900 2307 99030
rect 2627 94900 2667 99030
rect 2267 94860 2667 94900
rect -2766 94520 -2366 94560
rect -2766 90390 -2726 94520
rect -2406 90390 -2366 94520
rect -2766 90350 -2366 90390
rect -2047 94520 -1647 94560
rect -2047 90390 -2007 94520
rect -1687 90390 -1647 94520
rect -2047 90350 -1647 90390
rect -1328 94520 -928 94560
rect -1328 90390 -1288 94520
rect -968 90390 -928 94520
rect -1328 90350 -928 90390
rect -609 94520 -209 94560
rect -609 90390 -569 94520
rect -249 90390 -209 94520
rect -609 90350 -209 90390
rect 110 94520 510 94560
rect 110 90390 150 94520
rect 470 90390 510 94520
rect 110 90350 510 90390
rect 829 94520 1229 94560
rect 829 90390 869 94520
rect 1189 90390 1229 94520
rect 829 90350 1229 90390
rect 1548 94520 1948 94560
rect 1548 90390 1588 94520
rect 1908 90390 1948 94520
rect 1548 90350 1948 90390
rect 2267 94520 2667 94560
rect 2267 90390 2307 94520
rect 2627 90390 2667 94520
rect 2267 90350 2667 90390
rect -2766 90010 -2366 90050
rect -2766 85880 -2726 90010
rect -2406 85880 -2366 90010
rect -2766 85840 -2366 85880
rect -2047 90010 -1647 90050
rect -2047 85880 -2007 90010
rect -1687 85880 -1647 90010
rect -2047 85840 -1647 85880
rect -1328 90010 -928 90050
rect -1328 85880 -1288 90010
rect -968 85880 -928 90010
rect -1328 85840 -928 85880
rect -609 90010 -209 90050
rect -609 85880 -569 90010
rect -249 85880 -209 90010
rect -609 85840 -209 85880
rect 110 90010 510 90050
rect 110 85880 150 90010
rect 470 85880 510 90010
rect 110 85840 510 85880
rect 829 90010 1229 90050
rect 829 85880 869 90010
rect 1189 85880 1229 90010
rect 829 85840 1229 85880
rect 1548 90010 1948 90050
rect 1548 85880 1588 90010
rect 1908 85880 1948 90010
rect 1548 85840 1948 85880
rect 2267 90010 2667 90050
rect 2267 85880 2307 90010
rect 2627 85880 2667 90010
rect 2267 85840 2667 85880
rect -2766 85500 -2366 85540
rect -2766 81370 -2726 85500
rect -2406 81370 -2366 85500
rect -2766 81330 -2366 81370
rect -2047 85500 -1647 85540
rect -2047 81370 -2007 85500
rect -1687 81370 -1647 85500
rect -2047 81330 -1647 81370
rect -1328 85500 -928 85540
rect -1328 81370 -1288 85500
rect -968 81370 -928 85500
rect -1328 81330 -928 81370
rect -609 85500 -209 85540
rect -609 81370 -569 85500
rect -249 81370 -209 85500
rect -609 81330 -209 81370
rect 110 85500 510 85540
rect 110 81370 150 85500
rect 470 81370 510 85500
rect 110 81330 510 81370
rect 829 85500 1229 85540
rect 829 81370 869 85500
rect 1189 81370 1229 85500
rect 829 81330 1229 81370
rect 1548 85500 1948 85540
rect 1548 81370 1588 85500
rect 1908 81370 1948 85500
rect 1548 81330 1948 81370
rect 2267 85500 2667 85540
rect 2267 81370 2307 85500
rect 2627 81370 2667 85500
rect 2267 81330 2667 81370
rect -2766 80990 -2366 81030
rect -2766 76860 -2726 80990
rect -2406 76860 -2366 80990
rect -2766 76820 -2366 76860
rect -2047 80990 -1647 81030
rect -2047 76860 -2007 80990
rect -1687 76860 -1647 80990
rect -2047 76820 -1647 76860
rect -1328 80990 -928 81030
rect -1328 76860 -1288 80990
rect -968 76860 -928 80990
rect -1328 76820 -928 76860
rect -609 80990 -209 81030
rect -609 76860 -569 80990
rect -249 76860 -209 80990
rect -609 76820 -209 76860
rect 110 80990 510 81030
rect 110 76860 150 80990
rect 470 76860 510 80990
rect 110 76820 510 76860
rect 829 80990 1229 81030
rect 829 76860 869 80990
rect 1189 76860 1229 80990
rect 829 76820 1229 76860
rect 1548 80990 1948 81030
rect 1548 76860 1588 80990
rect 1908 76860 1948 80990
rect 1548 76820 1948 76860
rect 2267 80990 2667 81030
rect 2267 76860 2307 80990
rect 2627 76860 2667 80990
rect 2267 76820 2667 76860
rect -2766 76480 -2366 76520
rect -2766 72350 -2726 76480
rect -2406 72350 -2366 76480
rect -2766 72310 -2366 72350
rect -2047 76480 -1647 76520
rect -2047 72350 -2007 76480
rect -1687 72350 -1647 76480
rect -2047 72310 -1647 72350
rect -1328 76480 -928 76520
rect -1328 72350 -1288 76480
rect -968 72350 -928 76480
rect -1328 72310 -928 72350
rect -609 76480 -209 76520
rect -609 72350 -569 76480
rect -249 72350 -209 76480
rect -609 72310 -209 72350
rect 110 76480 510 76520
rect 110 72350 150 76480
rect 470 72350 510 76480
rect 110 72310 510 72350
rect 829 76480 1229 76520
rect 829 72350 869 76480
rect 1189 72350 1229 76480
rect 829 72310 1229 72350
rect 1548 76480 1948 76520
rect 1548 72350 1588 76480
rect 1908 72350 1948 76480
rect 1548 72310 1948 72350
rect 2267 76480 2667 76520
rect 2267 72350 2307 76480
rect 2627 72350 2667 76480
rect 2267 72310 2667 72350
rect -2766 71970 -2366 72010
rect -2766 67840 -2726 71970
rect -2406 67840 -2366 71970
rect -2766 67800 -2366 67840
rect -2047 71970 -1647 72010
rect -2047 67840 -2007 71970
rect -1687 67840 -1647 71970
rect -2047 67800 -1647 67840
rect -1328 71970 -928 72010
rect -1328 67840 -1288 71970
rect -968 67840 -928 71970
rect -1328 67800 -928 67840
rect -609 71970 -209 72010
rect -609 67840 -569 71970
rect -249 67840 -209 71970
rect -609 67800 -209 67840
rect 110 71970 510 72010
rect 110 67840 150 71970
rect 470 67840 510 71970
rect 110 67800 510 67840
rect 829 71970 1229 72010
rect 829 67840 869 71970
rect 1189 67840 1229 71970
rect 829 67800 1229 67840
rect 1548 71970 1948 72010
rect 1548 67840 1588 71970
rect 1908 67840 1948 71970
rect 1548 67800 1948 67840
rect 2267 71970 2667 72010
rect 2267 67840 2307 71970
rect 2627 67840 2667 71970
rect 2267 67800 2667 67840
rect -2766 67460 -2366 67500
rect -2766 63330 -2726 67460
rect -2406 63330 -2366 67460
rect -2766 63290 -2366 63330
rect -2047 67460 -1647 67500
rect -2047 63330 -2007 67460
rect -1687 63330 -1647 67460
rect -2047 63290 -1647 63330
rect -1328 67460 -928 67500
rect -1328 63330 -1288 67460
rect -968 63330 -928 67460
rect -1328 63290 -928 63330
rect -609 67460 -209 67500
rect -609 63330 -569 67460
rect -249 63330 -209 67460
rect -609 63290 -209 63330
rect 110 67460 510 67500
rect 110 63330 150 67460
rect 470 63330 510 67460
rect 110 63290 510 63330
rect 829 67460 1229 67500
rect 829 63330 869 67460
rect 1189 63330 1229 67460
rect 829 63290 1229 63330
rect 1548 67460 1948 67500
rect 1548 63330 1588 67460
rect 1908 63330 1948 67460
rect 1548 63290 1948 63330
rect 2267 67460 2667 67500
rect 2267 63330 2307 67460
rect 2627 63330 2667 67460
rect 2267 63290 2667 63330
rect -2766 62950 -2366 62990
rect -2766 58820 -2726 62950
rect -2406 58820 -2366 62950
rect -2766 58780 -2366 58820
rect -2047 62950 -1647 62990
rect -2047 58820 -2007 62950
rect -1687 58820 -1647 62950
rect -2047 58780 -1647 58820
rect -1328 62950 -928 62990
rect -1328 58820 -1288 62950
rect -968 58820 -928 62950
rect -1328 58780 -928 58820
rect -609 62950 -209 62990
rect -609 58820 -569 62950
rect -249 58820 -209 62950
rect -609 58780 -209 58820
rect 110 62950 510 62990
rect 110 58820 150 62950
rect 470 58820 510 62950
rect 110 58780 510 58820
rect 829 62950 1229 62990
rect 829 58820 869 62950
rect 1189 58820 1229 62950
rect 829 58780 1229 58820
rect 1548 62950 1948 62990
rect 1548 58820 1588 62950
rect 1908 58820 1948 62950
rect 1548 58780 1948 58820
rect 2267 62950 2667 62990
rect 2267 58820 2307 62950
rect 2627 58820 2667 62950
rect 2267 58780 2667 58820
rect -2766 58440 -2366 58480
rect -2766 54310 -2726 58440
rect -2406 54310 -2366 58440
rect -2766 54270 -2366 54310
rect -2047 58440 -1647 58480
rect -2047 54310 -2007 58440
rect -1687 54310 -1647 58440
rect -2047 54270 -1647 54310
rect -1328 58440 -928 58480
rect -1328 54310 -1288 58440
rect -968 54310 -928 58440
rect -1328 54270 -928 54310
rect -609 58440 -209 58480
rect -609 54310 -569 58440
rect -249 54310 -209 58440
rect -609 54270 -209 54310
rect 110 58440 510 58480
rect 110 54310 150 58440
rect 470 54310 510 58440
rect 110 54270 510 54310
rect 829 58440 1229 58480
rect 829 54310 869 58440
rect 1189 54310 1229 58440
rect 829 54270 1229 54310
rect 1548 58440 1948 58480
rect 1548 54310 1588 58440
rect 1908 54310 1948 58440
rect 1548 54270 1948 54310
rect 2267 58440 2667 58480
rect 2267 54310 2307 58440
rect 2627 54310 2667 58440
rect 2267 54270 2667 54310
rect -2766 53930 -2366 53970
rect -2766 49800 -2726 53930
rect -2406 49800 -2366 53930
rect -2766 49760 -2366 49800
rect -2047 53930 -1647 53970
rect -2047 49800 -2007 53930
rect -1687 49800 -1647 53930
rect -2047 49760 -1647 49800
rect -1328 53930 -928 53970
rect -1328 49800 -1288 53930
rect -968 49800 -928 53930
rect -1328 49760 -928 49800
rect -609 53930 -209 53970
rect -609 49800 -569 53930
rect -249 49800 -209 53930
rect -609 49760 -209 49800
rect 110 53930 510 53970
rect 110 49800 150 53930
rect 470 49800 510 53930
rect 110 49760 510 49800
rect 829 53930 1229 53970
rect 829 49800 869 53930
rect 1189 49800 1229 53930
rect 829 49760 1229 49800
rect 1548 53930 1948 53970
rect 1548 49800 1588 53930
rect 1908 49800 1948 53930
rect 1548 49760 1948 49800
rect 2267 53930 2667 53970
rect 2267 49800 2307 53930
rect 2627 49800 2667 53930
rect 2267 49760 2667 49800
rect -2766 49420 -2366 49460
rect -2766 45290 -2726 49420
rect -2406 45290 -2366 49420
rect -2766 45250 -2366 45290
rect -2047 49420 -1647 49460
rect -2047 45290 -2007 49420
rect -1687 45290 -1647 49420
rect -2047 45250 -1647 45290
rect -1328 49420 -928 49460
rect -1328 45290 -1288 49420
rect -968 45290 -928 49420
rect -1328 45250 -928 45290
rect -609 49420 -209 49460
rect -609 45290 -569 49420
rect -249 45290 -209 49420
rect -609 45250 -209 45290
rect 110 49420 510 49460
rect 110 45290 150 49420
rect 470 45290 510 49420
rect 110 45250 510 45290
rect 829 49420 1229 49460
rect 829 45290 869 49420
rect 1189 45290 1229 49420
rect 829 45250 1229 45290
rect 1548 49420 1948 49460
rect 1548 45290 1588 49420
rect 1908 45290 1948 49420
rect 1548 45250 1948 45290
rect 2267 49420 2667 49460
rect 2267 45290 2307 49420
rect 2627 45290 2667 49420
rect 2267 45250 2667 45290
rect -2766 44910 -2366 44950
rect -2766 40780 -2726 44910
rect -2406 40780 -2366 44910
rect -2766 40740 -2366 40780
rect -2047 44910 -1647 44950
rect -2047 40780 -2007 44910
rect -1687 40780 -1647 44910
rect -2047 40740 -1647 40780
rect -1328 44910 -928 44950
rect -1328 40780 -1288 44910
rect -968 40780 -928 44910
rect -1328 40740 -928 40780
rect -609 44910 -209 44950
rect -609 40780 -569 44910
rect -249 40780 -209 44910
rect -609 40740 -209 40780
rect 110 44910 510 44950
rect 110 40780 150 44910
rect 470 40780 510 44910
rect 110 40740 510 40780
rect 829 44910 1229 44950
rect 829 40780 869 44910
rect 1189 40780 1229 44910
rect 829 40740 1229 40780
rect 1548 44910 1948 44950
rect 1548 40780 1588 44910
rect 1908 40780 1948 44910
rect 1548 40740 1948 40780
rect 2267 44910 2667 44950
rect 2267 40780 2307 44910
rect 2627 40780 2667 44910
rect 2267 40740 2667 40780
rect -2766 40400 -2366 40440
rect -2766 36270 -2726 40400
rect -2406 36270 -2366 40400
rect -2766 36230 -2366 36270
rect -2047 40400 -1647 40440
rect -2047 36270 -2007 40400
rect -1687 36270 -1647 40400
rect -2047 36230 -1647 36270
rect -1328 40400 -928 40440
rect -1328 36270 -1288 40400
rect -968 36270 -928 40400
rect -1328 36230 -928 36270
rect -609 40400 -209 40440
rect -609 36270 -569 40400
rect -249 36270 -209 40400
rect -609 36230 -209 36270
rect 110 40400 510 40440
rect 110 36270 150 40400
rect 470 36270 510 40400
rect 110 36230 510 36270
rect 829 40400 1229 40440
rect 829 36270 869 40400
rect 1189 36270 1229 40400
rect 829 36230 1229 36270
rect 1548 40400 1948 40440
rect 1548 36270 1588 40400
rect 1908 36270 1948 40400
rect 1548 36230 1948 36270
rect 2267 40400 2667 40440
rect 2267 36270 2307 40400
rect 2627 36270 2667 40400
rect 2267 36230 2667 36270
rect -2766 35890 -2366 35930
rect -2766 31760 -2726 35890
rect -2406 31760 -2366 35890
rect -2766 31720 -2366 31760
rect -2047 35890 -1647 35930
rect -2047 31760 -2007 35890
rect -1687 31760 -1647 35890
rect -2047 31720 -1647 31760
rect -1328 35890 -928 35930
rect -1328 31760 -1288 35890
rect -968 31760 -928 35890
rect -1328 31720 -928 31760
rect -609 35890 -209 35930
rect -609 31760 -569 35890
rect -249 31760 -209 35890
rect -609 31720 -209 31760
rect 110 35890 510 35930
rect 110 31760 150 35890
rect 470 31760 510 35890
rect 110 31720 510 31760
rect 829 35890 1229 35930
rect 829 31760 869 35890
rect 1189 31760 1229 35890
rect 829 31720 1229 31760
rect 1548 35890 1948 35930
rect 1548 31760 1588 35890
rect 1908 31760 1948 35890
rect 1548 31720 1948 31760
rect 2267 35890 2667 35930
rect 2267 31760 2307 35890
rect 2627 31760 2667 35890
rect 2267 31720 2667 31760
rect -2766 31380 -2366 31420
rect -2766 27250 -2726 31380
rect -2406 27250 -2366 31380
rect -2766 27210 -2366 27250
rect -2047 31380 -1647 31420
rect -2047 27250 -2007 31380
rect -1687 27250 -1647 31380
rect -2047 27210 -1647 27250
rect -1328 31380 -928 31420
rect -1328 27250 -1288 31380
rect -968 27250 -928 31380
rect -1328 27210 -928 27250
rect -609 31380 -209 31420
rect -609 27250 -569 31380
rect -249 27250 -209 31380
rect -609 27210 -209 27250
rect 110 31380 510 31420
rect 110 27250 150 31380
rect 470 27250 510 31380
rect 110 27210 510 27250
rect 829 31380 1229 31420
rect 829 27250 869 31380
rect 1189 27250 1229 31380
rect 829 27210 1229 27250
rect 1548 31380 1948 31420
rect 1548 27250 1588 31380
rect 1908 27250 1948 31380
rect 1548 27210 1948 27250
rect 2267 31380 2667 31420
rect 2267 27250 2307 31380
rect 2627 27250 2667 31380
rect 2267 27210 2667 27250
rect -2766 26870 -2366 26910
rect -2766 22740 -2726 26870
rect -2406 22740 -2366 26870
rect -2766 22700 -2366 22740
rect -2047 26870 -1647 26910
rect -2047 22740 -2007 26870
rect -1687 22740 -1647 26870
rect -2047 22700 -1647 22740
rect -1328 26870 -928 26910
rect -1328 22740 -1288 26870
rect -968 22740 -928 26870
rect -1328 22700 -928 22740
rect -609 26870 -209 26910
rect -609 22740 -569 26870
rect -249 22740 -209 26870
rect -609 22700 -209 22740
rect 110 26870 510 26910
rect 110 22740 150 26870
rect 470 22740 510 26870
rect 110 22700 510 22740
rect 829 26870 1229 26910
rect 829 22740 869 26870
rect 1189 22740 1229 26870
rect 829 22700 1229 22740
rect 1548 26870 1948 26910
rect 1548 22740 1588 26870
rect 1908 22740 1948 26870
rect 1548 22700 1948 22740
rect 2267 26870 2667 26910
rect 2267 22740 2307 26870
rect 2627 22740 2667 26870
rect 2267 22700 2667 22740
rect -2766 22360 -2366 22400
rect -2766 18230 -2726 22360
rect -2406 18230 -2366 22360
rect -2766 18190 -2366 18230
rect -2047 22360 -1647 22400
rect -2047 18230 -2007 22360
rect -1687 18230 -1647 22360
rect -2047 18190 -1647 18230
rect -1328 22360 -928 22400
rect -1328 18230 -1288 22360
rect -968 18230 -928 22360
rect -1328 18190 -928 18230
rect -609 22360 -209 22400
rect -609 18230 -569 22360
rect -249 18230 -209 22360
rect -609 18190 -209 18230
rect 110 22360 510 22400
rect 110 18230 150 22360
rect 470 18230 510 22360
rect 110 18190 510 18230
rect 829 22360 1229 22400
rect 829 18230 869 22360
rect 1189 18230 1229 22360
rect 829 18190 1229 18230
rect 1548 22360 1948 22400
rect 1548 18230 1588 22360
rect 1908 18230 1948 22360
rect 1548 18190 1948 18230
rect 2267 22360 2667 22400
rect 2267 18230 2307 22360
rect 2627 18230 2667 22360
rect 2267 18190 2667 18230
rect -2766 17850 -2366 17890
rect -2766 13720 -2726 17850
rect -2406 13720 -2366 17850
rect -2766 13680 -2366 13720
rect -2047 17850 -1647 17890
rect -2047 13720 -2007 17850
rect -1687 13720 -1647 17850
rect -2047 13680 -1647 13720
rect -1328 17850 -928 17890
rect -1328 13720 -1288 17850
rect -968 13720 -928 17850
rect -1328 13680 -928 13720
rect -609 17850 -209 17890
rect -609 13720 -569 17850
rect -249 13720 -209 17850
rect -609 13680 -209 13720
rect 110 17850 510 17890
rect 110 13720 150 17850
rect 470 13720 510 17850
rect 110 13680 510 13720
rect 829 17850 1229 17890
rect 829 13720 869 17850
rect 1189 13720 1229 17850
rect 829 13680 1229 13720
rect 1548 17850 1948 17890
rect 1548 13720 1588 17850
rect 1908 13720 1948 17850
rect 1548 13680 1948 13720
rect 2267 17850 2667 17890
rect 2267 13720 2307 17850
rect 2627 13720 2667 17850
rect 2267 13680 2667 13720
rect -2766 13340 -2366 13380
rect -2766 9210 -2726 13340
rect -2406 9210 -2366 13340
rect -2766 9170 -2366 9210
rect -2047 13340 -1647 13380
rect -2047 9210 -2007 13340
rect -1687 9210 -1647 13340
rect -2047 9170 -1647 9210
rect -1328 13340 -928 13380
rect -1328 9210 -1288 13340
rect -968 9210 -928 13340
rect -1328 9170 -928 9210
rect -609 13340 -209 13380
rect -609 9210 -569 13340
rect -249 9210 -209 13340
rect -609 9170 -209 9210
rect 110 13340 510 13380
rect 110 9210 150 13340
rect 470 9210 510 13340
rect 110 9170 510 9210
rect 829 13340 1229 13380
rect 829 9210 869 13340
rect 1189 9210 1229 13340
rect 829 9170 1229 9210
rect 1548 13340 1948 13380
rect 1548 9210 1588 13340
rect 1908 9210 1948 13340
rect 1548 9170 1948 9210
rect 2267 13340 2667 13380
rect 2267 9210 2307 13340
rect 2627 9210 2667 13340
rect 2267 9170 2667 9210
rect -2766 8830 -2366 8870
rect -2766 4700 -2726 8830
rect -2406 4700 -2366 8830
rect -2766 4660 -2366 4700
rect -2047 8830 -1647 8870
rect -2047 4700 -2007 8830
rect -1687 4700 -1647 8830
rect -2047 4660 -1647 4700
rect -1328 8830 -928 8870
rect -1328 4700 -1288 8830
rect -968 4700 -928 8830
rect -1328 4660 -928 4700
rect -609 8830 -209 8870
rect -609 4700 -569 8830
rect -249 4700 -209 8830
rect -609 4660 -209 4700
rect 110 8830 510 8870
rect 110 4700 150 8830
rect 470 4700 510 8830
rect 110 4660 510 4700
rect 829 8830 1229 8870
rect 829 4700 869 8830
rect 1189 4700 1229 8830
rect 829 4660 1229 4700
rect 1548 8830 1948 8870
rect 1548 4700 1588 8830
rect 1908 4700 1948 8830
rect 1548 4660 1948 4700
rect 2267 8830 2667 8870
rect 2267 4700 2307 8830
rect 2627 4700 2667 8830
rect 2267 4660 2667 4700
rect -2766 4320 -2366 4360
rect -2766 190 -2726 4320
rect -2406 190 -2366 4320
rect -2766 150 -2366 190
rect -2047 4320 -1647 4360
rect -2047 190 -2007 4320
rect -1687 190 -1647 4320
rect -2047 150 -1647 190
rect -1328 4320 -928 4360
rect -1328 190 -1288 4320
rect -968 190 -928 4320
rect -1328 150 -928 190
rect -609 4320 -209 4360
rect -609 190 -569 4320
rect -249 190 -209 4320
rect -609 150 -209 190
rect 110 4320 510 4360
rect 110 190 150 4320
rect 470 190 510 4320
rect 110 150 510 190
rect 829 4320 1229 4360
rect 829 190 869 4320
rect 1189 190 1229 4320
rect 829 150 1229 190
rect 1548 4320 1948 4360
rect 1548 190 1588 4320
rect 1908 190 1948 4320
rect 1548 150 1948 190
rect 2267 4320 2667 4360
rect 2267 190 2307 4320
rect 2627 190 2667 4320
rect 2267 150 2667 190
rect -2766 -190 -2366 -150
rect -2766 -4320 -2726 -190
rect -2406 -4320 -2366 -190
rect -2766 -4360 -2366 -4320
rect -2047 -190 -1647 -150
rect -2047 -4320 -2007 -190
rect -1687 -4320 -1647 -190
rect -2047 -4360 -1647 -4320
rect -1328 -190 -928 -150
rect -1328 -4320 -1288 -190
rect -968 -4320 -928 -190
rect -1328 -4360 -928 -4320
rect -609 -190 -209 -150
rect -609 -4320 -569 -190
rect -249 -4320 -209 -190
rect -609 -4360 -209 -4320
rect 110 -190 510 -150
rect 110 -4320 150 -190
rect 470 -4320 510 -190
rect 110 -4360 510 -4320
rect 829 -190 1229 -150
rect 829 -4320 869 -190
rect 1189 -4320 1229 -190
rect 829 -4360 1229 -4320
rect 1548 -190 1948 -150
rect 1548 -4320 1588 -190
rect 1908 -4320 1948 -190
rect 1548 -4360 1948 -4320
rect 2267 -190 2667 -150
rect 2267 -4320 2307 -190
rect 2627 -4320 2667 -190
rect 2267 -4360 2667 -4320
rect -2766 -4700 -2366 -4660
rect -2766 -8830 -2726 -4700
rect -2406 -8830 -2366 -4700
rect -2766 -8870 -2366 -8830
rect -2047 -4700 -1647 -4660
rect -2047 -8830 -2007 -4700
rect -1687 -8830 -1647 -4700
rect -2047 -8870 -1647 -8830
rect -1328 -4700 -928 -4660
rect -1328 -8830 -1288 -4700
rect -968 -8830 -928 -4700
rect -1328 -8870 -928 -8830
rect -609 -4700 -209 -4660
rect -609 -8830 -569 -4700
rect -249 -8830 -209 -4700
rect -609 -8870 -209 -8830
rect 110 -4700 510 -4660
rect 110 -8830 150 -4700
rect 470 -8830 510 -4700
rect 110 -8870 510 -8830
rect 829 -4700 1229 -4660
rect 829 -8830 869 -4700
rect 1189 -8830 1229 -4700
rect 829 -8870 1229 -8830
rect 1548 -4700 1948 -4660
rect 1548 -8830 1588 -4700
rect 1908 -8830 1948 -4700
rect 1548 -8870 1948 -8830
rect 2267 -4700 2667 -4660
rect 2267 -8830 2307 -4700
rect 2627 -8830 2667 -4700
rect 2267 -8870 2667 -8830
rect -2766 -9210 -2366 -9170
rect -2766 -13340 -2726 -9210
rect -2406 -13340 -2366 -9210
rect -2766 -13380 -2366 -13340
rect -2047 -9210 -1647 -9170
rect -2047 -13340 -2007 -9210
rect -1687 -13340 -1647 -9210
rect -2047 -13380 -1647 -13340
rect -1328 -9210 -928 -9170
rect -1328 -13340 -1288 -9210
rect -968 -13340 -928 -9210
rect -1328 -13380 -928 -13340
rect -609 -9210 -209 -9170
rect -609 -13340 -569 -9210
rect -249 -13340 -209 -9210
rect -609 -13380 -209 -13340
rect 110 -9210 510 -9170
rect 110 -13340 150 -9210
rect 470 -13340 510 -9210
rect 110 -13380 510 -13340
rect 829 -9210 1229 -9170
rect 829 -13340 869 -9210
rect 1189 -13340 1229 -9210
rect 829 -13380 1229 -13340
rect 1548 -9210 1948 -9170
rect 1548 -13340 1588 -9210
rect 1908 -13340 1948 -9210
rect 1548 -13380 1948 -13340
rect 2267 -9210 2667 -9170
rect 2267 -13340 2307 -9210
rect 2627 -13340 2667 -9210
rect 2267 -13380 2667 -13340
rect -2766 -13720 -2366 -13680
rect -2766 -17850 -2726 -13720
rect -2406 -17850 -2366 -13720
rect -2766 -17890 -2366 -17850
rect -2047 -13720 -1647 -13680
rect -2047 -17850 -2007 -13720
rect -1687 -17850 -1647 -13720
rect -2047 -17890 -1647 -17850
rect -1328 -13720 -928 -13680
rect -1328 -17850 -1288 -13720
rect -968 -17850 -928 -13720
rect -1328 -17890 -928 -17850
rect -609 -13720 -209 -13680
rect -609 -17850 -569 -13720
rect -249 -17850 -209 -13720
rect -609 -17890 -209 -17850
rect 110 -13720 510 -13680
rect 110 -17850 150 -13720
rect 470 -17850 510 -13720
rect 110 -17890 510 -17850
rect 829 -13720 1229 -13680
rect 829 -17850 869 -13720
rect 1189 -17850 1229 -13720
rect 829 -17890 1229 -17850
rect 1548 -13720 1948 -13680
rect 1548 -17850 1588 -13720
rect 1908 -17850 1948 -13720
rect 1548 -17890 1948 -17850
rect 2267 -13720 2667 -13680
rect 2267 -17850 2307 -13720
rect 2627 -17850 2667 -13720
rect 2267 -17890 2667 -17850
rect -2766 -18230 -2366 -18190
rect -2766 -22360 -2726 -18230
rect -2406 -22360 -2366 -18230
rect -2766 -22400 -2366 -22360
rect -2047 -18230 -1647 -18190
rect -2047 -22360 -2007 -18230
rect -1687 -22360 -1647 -18230
rect -2047 -22400 -1647 -22360
rect -1328 -18230 -928 -18190
rect -1328 -22360 -1288 -18230
rect -968 -22360 -928 -18230
rect -1328 -22400 -928 -22360
rect -609 -18230 -209 -18190
rect -609 -22360 -569 -18230
rect -249 -22360 -209 -18230
rect -609 -22400 -209 -22360
rect 110 -18230 510 -18190
rect 110 -22360 150 -18230
rect 470 -22360 510 -18230
rect 110 -22400 510 -22360
rect 829 -18230 1229 -18190
rect 829 -22360 869 -18230
rect 1189 -22360 1229 -18230
rect 829 -22400 1229 -22360
rect 1548 -18230 1948 -18190
rect 1548 -22360 1588 -18230
rect 1908 -22360 1948 -18230
rect 1548 -22400 1948 -22360
rect 2267 -18230 2667 -18190
rect 2267 -22360 2307 -18230
rect 2627 -22360 2667 -18230
rect 2267 -22400 2667 -22360
rect -2766 -22740 -2366 -22700
rect -2766 -26870 -2726 -22740
rect -2406 -26870 -2366 -22740
rect -2766 -26910 -2366 -26870
rect -2047 -22740 -1647 -22700
rect -2047 -26870 -2007 -22740
rect -1687 -26870 -1647 -22740
rect -2047 -26910 -1647 -26870
rect -1328 -22740 -928 -22700
rect -1328 -26870 -1288 -22740
rect -968 -26870 -928 -22740
rect -1328 -26910 -928 -26870
rect -609 -22740 -209 -22700
rect -609 -26870 -569 -22740
rect -249 -26870 -209 -22740
rect -609 -26910 -209 -26870
rect 110 -22740 510 -22700
rect 110 -26870 150 -22740
rect 470 -26870 510 -22740
rect 110 -26910 510 -26870
rect 829 -22740 1229 -22700
rect 829 -26870 869 -22740
rect 1189 -26870 1229 -22740
rect 829 -26910 1229 -26870
rect 1548 -22740 1948 -22700
rect 1548 -26870 1588 -22740
rect 1908 -26870 1948 -22740
rect 1548 -26910 1948 -26870
rect 2267 -22740 2667 -22700
rect 2267 -26870 2307 -22740
rect 2627 -26870 2667 -22740
rect 2267 -26910 2667 -26870
rect -2766 -27250 -2366 -27210
rect -2766 -31380 -2726 -27250
rect -2406 -31380 -2366 -27250
rect -2766 -31420 -2366 -31380
rect -2047 -27250 -1647 -27210
rect -2047 -31380 -2007 -27250
rect -1687 -31380 -1647 -27250
rect -2047 -31420 -1647 -31380
rect -1328 -27250 -928 -27210
rect -1328 -31380 -1288 -27250
rect -968 -31380 -928 -27250
rect -1328 -31420 -928 -31380
rect -609 -27250 -209 -27210
rect -609 -31380 -569 -27250
rect -249 -31380 -209 -27250
rect -609 -31420 -209 -31380
rect 110 -27250 510 -27210
rect 110 -31380 150 -27250
rect 470 -31380 510 -27250
rect 110 -31420 510 -31380
rect 829 -27250 1229 -27210
rect 829 -31380 869 -27250
rect 1189 -31380 1229 -27250
rect 829 -31420 1229 -31380
rect 1548 -27250 1948 -27210
rect 1548 -31380 1588 -27250
rect 1908 -31380 1948 -27250
rect 1548 -31420 1948 -31380
rect 2267 -27250 2667 -27210
rect 2267 -31380 2307 -27250
rect 2627 -31380 2667 -27250
rect 2267 -31420 2667 -31380
rect -2766 -31760 -2366 -31720
rect -2766 -35890 -2726 -31760
rect -2406 -35890 -2366 -31760
rect -2766 -35930 -2366 -35890
rect -2047 -31760 -1647 -31720
rect -2047 -35890 -2007 -31760
rect -1687 -35890 -1647 -31760
rect -2047 -35930 -1647 -35890
rect -1328 -31760 -928 -31720
rect -1328 -35890 -1288 -31760
rect -968 -35890 -928 -31760
rect -1328 -35930 -928 -35890
rect -609 -31760 -209 -31720
rect -609 -35890 -569 -31760
rect -249 -35890 -209 -31760
rect -609 -35930 -209 -35890
rect 110 -31760 510 -31720
rect 110 -35890 150 -31760
rect 470 -35890 510 -31760
rect 110 -35930 510 -35890
rect 829 -31760 1229 -31720
rect 829 -35890 869 -31760
rect 1189 -35890 1229 -31760
rect 829 -35930 1229 -35890
rect 1548 -31760 1948 -31720
rect 1548 -35890 1588 -31760
rect 1908 -35890 1948 -31760
rect 1548 -35930 1948 -35890
rect 2267 -31760 2667 -31720
rect 2267 -35890 2307 -31760
rect 2627 -35890 2667 -31760
rect 2267 -35930 2667 -35890
rect -2766 -36270 -2366 -36230
rect -2766 -40400 -2726 -36270
rect -2406 -40400 -2366 -36270
rect -2766 -40440 -2366 -40400
rect -2047 -36270 -1647 -36230
rect -2047 -40400 -2007 -36270
rect -1687 -40400 -1647 -36270
rect -2047 -40440 -1647 -40400
rect -1328 -36270 -928 -36230
rect -1328 -40400 -1288 -36270
rect -968 -40400 -928 -36270
rect -1328 -40440 -928 -40400
rect -609 -36270 -209 -36230
rect -609 -40400 -569 -36270
rect -249 -40400 -209 -36270
rect -609 -40440 -209 -40400
rect 110 -36270 510 -36230
rect 110 -40400 150 -36270
rect 470 -40400 510 -36270
rect 110 -40440 510 -40400
rect 829 -36270 1229 -36230
rect 829 -40400 869 -36270
rect 1189 -40400 1229 -36270
rect 829 -40440 1229 -40400
rect 1548 -36270 1948 -36230
rect 1548 -40400 1588 -36270
rect 1908 -40400 1948 -36270
rect 1548 -40440 1948 -40400
rect 2267 -36270 2667 -36230
rect 2267 -40400 2307 -36270
rect 2627 -40400 2667 -36270
rect 2267 -40440 2667 -40400
rect -2766 -40780 -2366 -40740
rect -2766 -44910 -2726 -40780
rect -2406 -44910 -2366 -40780
rect -2766 -44950 -2366 -44910
rect -2047 -40780 -1647 -40740
rect -2047 -44910 -2007 -40780
rect -1687 -44910 -1647 -40780
rect -2047 -44950 -1647 -44910
rect -1328 -40780 -928 -40740
rect -1328 -44910 -1288 -40780
rect -968 -44910 -928 -40780
rect -1328 -44950 -928 -44910
rect -609 -40780 -209 -40740
rect -609 -44910 -569 -40780
rect -249 -44910 -209 -40780
rect -609 -44950 -209 -44910
rect 110 -40780 510 -40740
rect 110 -44910 150 -40780
rect 470 -44910 510 -40780
rect 110 -44950 510 -44910
rect 829 -40780 1229 -40740
rect 829 -44910 869 -40780
rect 1189 -44910 1229 -40780
rect 829 -44950 1229 -44910
rect 1548 -40780 1948 -40740
rect 1548 -44910 1588 -40780
rect 1908 -44910 1948 -40780
rect 1548 -44950 1948 -44910
rect 2267 -40780 2667 -40740
rect 2267 -44910 2307 -40780
rect 2627 -44910 2667 -40780
rect 2267 -44950 2667 -44910
rect -2766 -45290 -2366 -45250
rect -2766 -49420 -2726 -45290
rect -2406 -49420 -2366 -45290
rect -2766 -49460 -2366 -49420
rect -2047 -45290 -1647 -45250
rect -2047 -49420 -2007 -45290
rect -1687 -49420 -1647 -45290
rect -2047 -49460 -1647 -49420
rect -1328 -45290 -928 -45250
rect -1328 -49420 -1288 -45290
rect -968 -49420 -928 -45290
rect -1328 -49460 -928 -49420
rect -609 -45290 -209 -45250
rect -609 -49420 -569 -45290
rect -249 -49420 -209 -45290
rect -609 -49460 -209 -49420
rect 110 -45290 510 -45250
rect 110 -49420 150 -45290
rect 470 -49420 510 -45290
rect 110 -49460 510 -49420
rect 829 -45290 1229 -45250
rect 829 -49420 869 -45290
rect 1189 -49420 1229 -45290
rect 829 -49460 1229 -49420
rect 1548 -45290 1948 -45250
rect 1548 -49420 1588 -45290
rect 1908 -49420 1948 -45290
rect 1548 -49460 1948 -49420
rect 2267 -45290 2667 -45250
rect 2267 -49420 2307 -45290
rect 2627 -49420 2667 -45290
rect 2267 -49460 2667 -49420
rect -2766 -49800 -2366 -49760
rect -2766 -53930 -2726 -49800
rect -2406 -53930 -2366 -49800
rect -2766 -53970 -2366 -53930
rect -2047 -49800 -1647 -49760
rect -2047 -53930 -2007 -49800
rect -1687 -53930 -1647 -49800
rect -2047 -53970 -1647 -53930
rect -1328 -49800 -928 -49760
rect -1328 -53930 -1288 -49800
rect -968 -53930 -928 -49800
rect -1328 -53970 -928 -53930
rect -609 -49800 -209 -49760
rect -609 -53930 -569 -49800
rect -249 -53930 -209 -49800
rect -609 -53970 -209 -53930
rect 110 -49800 510 -49760
rect 110 -53930 150 -49800
rect 470 -53930 510 -49800
rect 110 -53970 510 -53930
rect 829 -49800 1229 -49760
rect 829 -53930 869 -49800
rect 1189 -53930 1229 -49800
rect 829 -53970 1229 -53930
rect 1548 -49800 1948 -49760
rect 1548 -53930 1588 -49800
rect 1908 -53930 1948 -49800
rect 1548 -53970 1948 -53930
rect 2267 -49800 2667 -49760
rect 2267 -53930 2307 -49800
rect 2627 -53930 2667 -49800
rect 2267 -53970 2667 -53930
rect -2766 -54310 -2366 -54270
rect -2766 -58440 -2726 -54310
rect -2406 -58440 -2366 -54310
rect -2766 -58480 -2366 -58440
rect -2047 -54310 -1647 -54270
rect -2047 -58440 -2007 -54310
rect -1687 -58440 -1647 -54310
rect -2047 -58480 -1647 -58440
rect -1328 -54310 -928 -54270
rect -1328 -58440 -1288 -54310
rect -968 -58440 -928 -54310
rect -1328 -58480 -928 -58440
rect -609 -54310 -209 -54270
rect -609 -58440 -569 -54310
rect -249 -58440 -209 -54310
rect -609 -58480 -209 -58440
rect 110 -54310 510 -54270
rect 110 -58440 150 -54310
rect 470 -58440 510 -54310
rect 110 -58480 510 -58440
rect 829 -54310 1229 -54270
rect 829 -58440 869 -54310
rect 1189 -58440 1229 -54310
rect 829 -58480 1229 -58440
rect 1548 -54310 1948 -54270
rect 1548 -58440 1588 -54310
rect 1908 -58440 1948 -54310
rect 1548 -58480 1948 -58440
rect 2267 -54310 2667 -54270
rect 2267 -58440 2307 -54310
rect 2627 -58440 2667 -54310
rect 2267 -58480 2667 -58440
rect -2766 -58820 -2366 -58780
rect -2766 -62950 -2726 -58820
rect -2406 -62950 -2366 -58820
rect -2766 -62990 -2366 -62950
rect -2047 -58820 -1647 -58780
rect -2047 -62950 -2007 -58820
rect -1687 -62950 -1647 -58820
rect -2047 -62990 -1647 -62950
rect -1328 -58820 -928 -58780
rect -1328 -62950 -1288 -58820
rect -968 -62950 -928 -58820
rect -1328 -62990 -928 -62950
rect -609 -58820 -209 -58780
rect -609 -62950 -569 -58820
rect -249 -62950 -209 -58820
rect -609 -62990 -209 -62950
rect 110 -58820 510 -58780
rect 110 -62950 150 -58820
rect 470 -62950 510 -58820
rect 110 -62990 510 -62950
rect 829 -58820 1229 -58780
rect 829 -62950 869 -58820
rect 1189 -62950 1229 -58820
rect 829 -62990 1229 -62950
rect 1548 -58820 1948 -58780
rect 1548 -62950 1588 -58820
rect 1908 -62950 1948 -58820
rect 1548 -62990 1948 -62950
rect 2267 -58820 2667 -58780
rect 2267 -62950 2307 -58820
rect 2627 -62950 2667 -58820
rect 2267 -62990 2667 -62950
rect -2766 -63330 -2366 -63290
rect -2766 -67460 -2726 -63330
rect -2406 -67460 -2366 -63330
rect -2766 -67500 -2366 -67460
rect -2047 -63330 -1647 -63290
rect -2047 -67460 -2007 -63330
rect -1687 -67460 -1647 -63330
rect -2047 -67500 -1647 -67460
rect -1328 -63330 -928 -63290
rect -1328 -67460 -1288 -63330
rect -968 -67460 -928 -63330
rect -1328 -67500 -928 -67460
rect -609 -63330 -209 -63290
rect -609 -67460 -569 -63330
rect -249 -67460 -209 -63330
rect -609 -67500 -209 -67460
rect 110 -63330 510 -63290
rect 110 -67460 150 -63330
rect 470 -67460 510 -63330
rect 110 -67500 510 -67460
rect 829 -63330 1229 -63290
rect 829 -67460 869 -63330
rect 1189 -67460 1229 -63330
rect 829 -67500 1229 -67460
rect 1548 -63330 1948 -63290
rect 1548 -67460 1588 -63330
rect 1908 -67460 1948 -63330
rect 1548 -67500 1948 -67460
rect 2267 -63330 2667 -63290
rect 2267 -67460 2307 -63330
rect 2627 -67460 2667 -63330
rect 2267 -67500 2667 -67460
rect -2766 -67840 -2366 -67800
rect -2766 -71970 -2726 -67840
rect -2406 -71970 -2366 -67840
rect -2766 -72010 -2366 -71970
rect -2047 -67840 -1647 -67800
rect -2047 -71970 -2007 -67840
rect -1687 -71970 -1647 -67840
rect -2047 -72010 -1647 -71970
rect -1328 -67840 -928 -67800
rect -1328 -71970 -1288 -67840
rect -968 -71970 -928 -67840
rect -1328 -72010 -928 -71970
rect -609 -67840 -209 -67800
rect -609 -71970 -569 -67840
rect -249 -71970 -209 -67840
rect -609 -72010 -209 -71970
rect 110 -67840 510 -67800
rect 110 -71970 150 -67840
rect 470 -71970 510 -67840
rect 110 -72010 510 -71970
rect 829 -67840 1229 -67800
rect 829 -71970 869 -67840
rect 1189 -71970 1229 -67840
rect 829 -72010 1229 -71970
rect 1548 -67840 1948 -67800
rect 1548 -71970 1588 -67840
rect 1908 -71970 1948 -67840
rect 1548 -72010 1948 -71970
rect 2267 -67840 2667 -67800
rect 2267 -71970 2307 -67840
rect 2627 -71970 2667 -67840
rect 2267 -72010 2667 -71970
rect -2766 -72350 -2366 -72310
rect -2766 -76480 -2726 -72350
rect -2406 -76480 -2366 -72350
rect -2766 -76520 -2366 -76480
rect -2047 -72350 -1647 -72310
rect -2047 -76480 -2007 -72350
rect -1687 -76480 -1647 -72350
rect -2047 -76520 -1647 -76480
rect -1328 -72350 -928 -72310
rect -1328 -76480 -1288 -72350
rect -968 -76480 -928 -72350
rect -1328 -76520 -928 -76480
rect -609 -72350 -209 -72310
rect -609 -76480 -569 -72350
rect -249 -76480 -209 -72350
rect -609 -76520 -209 -76480
rect 110 -72350 510 -72310
rect 110 -76480 150 -72350
rect 470 -76480 510 -72350
rect 110 -76520 510 -76480
rect 829 -72350 1229 -72310
rect 829 -76480 869 -72350
rect 1189 -76480 1229 -72350
rect 829 -76520 1229 -76480
rect 1548 -72350 1948 -72310
rect 1548 -76480 1588 -72350
rect 1908 -76480 1948 -72350
rect 1548 -76520 1948 -76480
rect 2267 -72350 2667 -72310
rect 2267 -76480 2307 -72350
rect 2627 -76480 2667 -72350
rect 2267 -76520 2667 -76480
rect -2766 -76860 -2366 -76820
rect -2766 -80990 -2726 -76860
rect -2406 -80990 -2366 -76860
rect -2766 -81030 -2366 -80990
rect -2047 -76860 -1647 -76820
rect -2047 -80990 -2007 -76860
rect -1687 -80990 -1647 -76860
rect -2047 -81030 -1647 -80990
rect -1328 -76860 -928 -76820
rect -1328 -80990 -1288 -76860
rect -968 -80990 -928 -76860
rect -1328 -81030 -928 -80990
rect -609 -76860 -209 -76820
rect -609 -80990 -569 -76860
rect -249 -80990 -209 -76860
rect -609 -81030 -209 -80990
rect 110 -76860 510 -76820
rect 110 -80990 150 -76860
rect 470 -80990 510 -76860
rect 110 -81030 510 -80990
rect 829 -76860 1229 -76820
rect 829 -80990 869 -76860
rect 1189 -80990 1229 -76860
rect 829 -81030 1229 -80990
rect 1548 -76860 1948 -76820
rect 1548 -80990 1588 -76860
rect 1908 -80990 1948 -76860
rect 1548 -81030 1948 -80990
rect 2267 -76860 2667 -76820
rect 2267 -80990 2307 -76860
rect 2627 -80990 2667 -76860
rect 2267 -81030 2667 -80990
rect -2766 -81370 -2366 -81330
rect -2766 -85500 -2726 -81370
rect -2406 -85500 -2366 -81370
rect -2766 -85540 -2366 -85500
rect -2047 -81370 -1647 -81330
rect -2047 -85500 -2007 -81370
rect -1687 -85500 -1647 -81370
rect -2047 -85540 -1647 -85500
rect -1328 -81370 -928 -81330
rect -1328 -85500 -1288 -81370
rect -968 -85500 -928 -81370
rect -1328 -85540 -928 -85500
rect -609 -81370 -209 -81330
rect -609 -85500 -569 -81370
rect -249 -85500 -209 -81370
rect -609 -85540 -209 -85500
rect 110 -81370 510 -81330
rect 110 -85500 150 -81370
rect 470 -85500 510 -81370
rect 110 -85540 510 -85500
rect 829 -81370 1229 -81330
rect 829 -85500 869 -81370
rect 1189 -85500 1229 -81370
rect 829 -85540 1229 -85500
rect 1548 -81370 1948 -81330
rect 1548 -85500 1588 -81370
rect 1908 -85500 1948 -81370
rect 1548 -85540 1948 -85500
rect 2267 -81370 2667 -81330
rect 2267 -85500 2307 -81370
rect 2627 -85500 2667 -81370
rect 2267 -85540 2667 -85500
rect -2766 -85880 -2366 -85840
rect -2766 -90010 -2726 -85880
rect -2406 -90010 -2366 -85880
rect -2766 -90050 -2366 -90010
rect -2047 -85880 -1647 -85840
rect -2047 -90010 -2007 -85880
rect -1687 -90010 -1647 -85880
rect -2047 -90050 -1647 -90010
rect -1328 -85880 -928 -85840
rect -1328 -90010 -1288 -85880
rect -968 -90010 -928 -85880
rect -1328 -90050 -928 -90010
rect -609 -85880 -209 -85840
rect -609 -90010 -569 -85880
rect -249 -90010 -209 -85880
rect -609 -90050 -209 -90010
rect 110 -85880 510 -85840
rect 110 -90010 150 -85880
rect 470 -90010 510 -85880
rect 110 -90050 510 -90010
rect 829 -85880 1229 -85840
rect 829 -90010 869 -85880
rect 1189 -90010 1229 -85880
rect 829 -90050 1229 -90010
rect 1548 -85880 1948 -85840
rect 1548 -90010 1588 -85880
rect 1908 -90010 1948 -85880
rect 1548 -90050 1948 -90010
rect 2267 -85880 2667 -85840
rect 2267 -90010 2307 -85880
rect 2627 -90010 2667 -85880
rect 2267 -90050 2667 -90010
rect -2766 -90390 -2366 -90350
rect -2766 -94520 -2726 -90390
rect -2406 -94520 -2366 -90390
rect -2766 -94560 -2366 -94520
rect -2047 -90390 -1647 -90350
rect -2047 -94520 -2007 -90390
rect -1687 -94520 -1647 -90390
rect -2047 -94560 -1647 -94520
rect -1328 -90390 -928 -90350
rect -1328 -94520 -1288 -90390
rect -968 -94520 -928 -90390
rect -1328 -94560 -928 -94520
rect -609 -90390 -209 -90350
rect -609 -94520 -569 -90390
rect -249 -94520 -209 -90390
rect -609 -94560 -209 -94520
rect 110 -90390 510 -90350
rect 110 -94520 150 -90390
rect 470 -94520 510 -90390
rect 110 -94560 510 -94520
rect 829 -90390 1229 -90350
rect 829 -94520 869 -90390
rect 1189 -94520 1229 -90390
rect 829 -94560 1229 -94520
rect 1548 -90390 1948 -90350
rect 1548 -94520 1588 -90390
rect 1908 -94520 1948 -90390
rect 1548 -94560 1948 -94520
rect 2267 -90390 2667 -90350
rect 2267 -94520 2307 -90390
rect 2627 -94520 2667 -90390
rect 2267 -94560 2667 -94520
rect -2766 -94900 -2366 -94860
rect -2766 -99030 -2726 -94900
rect -2406 -99030 -2366 -94900
rect -2766 -99070 -2366 -99030
rect -2047 -94900 -1647 -94860
rect -2047 -99030 -2007 -94900
rect -1687 -99030 -1647 -94900
rect -2047 -99070 -1647 -99030
rect -1328 -94900 -928 -94860
rect -1328 -99030 -1288 -94900
rect -968 -99030 -928 -94900
rect -1328 -99070 -928 -99030
rect -609 -94900 -209 -94860
rect -609 -99030 -569 -94900
rect -249 -99030 -209 -94900
rect -609 -99070 -209 -99030
rect 110 -94900 510 -94860
rect 110 -99030 150 -94900
rect 470 -99030 510 -94900
rect 110 -99070 510 -99030
rect 829 -94900 1229 -94860
rect 829 -99030 869 -94900
rect 1189 -99030 1229 -94900
rect 829 -99070 1229 -99030
rect 1548 -94900 1948 -94860
rect 1548 -99030 1588 -94900
rect 1908 -99030 1948 -94900
rect 1548 -99070 1948 -99030
rect 2267 -94900 2667 -94860
rect 2267 -99030 2307 -94900
rect 2627 -99030 2667 -94900
rect 2267 -99070 2667 -99030
rect -2766 -99410 -2366 -99370
rect -2766 -103540 -2726 -99410
rect -2406 -103540 -2366 -99410
rect -2766 -103580 -2366 -103540
rect -2047 -99410 -1647 -99370
rect -2047 -103540 -2007 -99410
rect -1687 -103540 -1647 -99410
rect -2047 -103580 -1647 -103540
rect -1328 -99410 -928 -99370
rect -1328 -103540 -1288 -99410
rect -968 -103540 -928 -99410
rect -1328 -103580 -928 -103540
rect -609 -99410 -209 -99370
rect -609 -103540 -569 -99410
rect -249 -103540 -209 -99410
rect -609 -103580 -209 -103540
rect 110 -99410 510 -99370
rect 110 -103540 150 -99410
rect 470 -103540 510 -99410
rect 110 -103580 510 -103540
rect 829 -99410 1229 -99370
rect 829 -103540 869 -99410
rect 1189 -103540 1229 -99410
rect 829 -103580 1229 -103540
rect 1548 -99410 1948 -99370
rect 1548 -103540 1588 -99410
rect 1908 -103540 1948 -99410
rect 1548 -103580 1948 -103540
rect 2267 -99410 2667 -99370
rect 2267 -103540 2307 -99410
rect 2627 -103540 2667 -99410
rect 2267 -103580 2667 -103540
rect -2766 -103920 -2366 -103880
rect -2766 -108050 -2726 -103920
rect -2406 -108050 -2366 -103920
rect -2766 -108090 -2366 -108050
rect -2047 -103920 -1647 -103880
rect -2047 -108050 -2007 -103920
rect -1687 -108050 -1647 -103920
rect -2047 -108090 -1647 -108050
rect -1328 -103920 -928 -103880
rect -1328 -108050 -1288 -103920
rect -968 -108050 -928 -103920
rect -1328 -108090 -928 -108050
rect -609 -103920 -209 -103880
rect -609 -108050 -569 -103920
rect -249 -108050 -209 -103920
rect -609 -108090 -209 -108050
rect 110 -103920 510 -103880
rect 110 -108050 150 -103920
rect 470 -108050 510 -103920
rect 110 -108090 510 -108050
rect 829 -103920 1229 -103880
rect 829 -108050 869 -103920
rect 1189 -108050 1229 -103920
rect 829 -108090 1229 -108050
rect 1548 -103920 1948 -103880
rect 1548 -108050 1588 -103920
rect 1908 -108050 1948 -103920
rect 1548 -108090 1948 -108050
rect 2267 -103920 2667 -103880
rect 2267 -108050 2307 -103920
rect 2627 -108050 2667 -103920
rect 2267 -108090 2667 -108050
rect -2766 -108430 -2366 -108390
rect -2766 -112560 -2726 -108430
rect -2406 -112560 -2366 -108430
rect -2766 -112600 -2366 -112560
rect -2047 -108430 -1647 -108390
rect -2047 -112560 -2007 -108430
rect -1687 -112560 -1647 -108430
rect -2047 -112600 -1647 -112560
rect -1328 -108430 -928 -108390
rect -1328 -112560 -1288 -108430
rect -968 -112560 -928 -108430
rect -1328 -112600 -928 -112560
rect -609 -108430 -209 -108390
rect -609 -112560 -569 -108430
rect -249 -112560 -209 -108430
rect -609 -112600 -209 -112560
rect 110 -108430 510 -108390
rect 110 -112560 150 -108430
rect 470 -112560 510 -108430
rect 110 -112600 510 -112560
rect 829 -108430 1229 -108390
rect 829 -112560 869 -108430
rect 1189 -112560 1229 -108430
rect 829 -112600 1229 -112560
rect 1548 -108430 1948 -108390
rect 1548 -112560 1588 -108430
rect 1908 -112560 1948 -108430
rect 1548 -112600 1948 -112560
rect 2267 -108430 2667 -108390
rect 2267 -112560 2307 -108430
rect 2627 -112560 2667 -108430
rect 2267 -112600 2667 -112560
rect -2766 -112940 -2366 -112900
rect -2766 -117070 -2726 -112940
rect -2406 -117070 -2366 -112940
rect -2766 -117110 -2366 -117070
rect -2047 -112940 -1647 -112900
rect -2047 -117070 -2007 -112940
rect -1687 -117070 -1647 -112940
rect -2047 -117110 -1647 -117070
rect -1328 -112940 -928 -112900
rect -1328 -117070 -1288 -112940
rect -968 -117070 -928 -112940
rect -1328 -117110 -928 -117070
rect -609 -112940 -209 -112900
rect -609 -117070 -569 -112940
rect -249 -117070 -209 -112940
rect -609 -117110 -209 -117070
rect 110 -112940 510 -112900
rect 110 -117070 150 -112940
rect 470 -117070 510 -112940
rect 110 -117110 510 -117070
rect 829 -112940 1229 -112900
rect 829 -117070 869 -112940
rect 1189 -117070 1229 -112940
rect 829 -117110 1229 -117070
rect 1548 -112940 1948 -112900
rect 1548 -117070 1588 -112940
rect 1908 -117070 1948 -112940
rect 1548 -117110 1948 -117070
rect 2267 -112940 2667 -112900
rect 2267 -117070 2307 -112940
rect 2627 -117070 2667 -112940
rect 2267 -117110 2667 -117070
rect -2766 -117450 -2366 -117410
rect -2766 -121580 -2726 -117450
rect -2406 -121580 -2366 -117450
rect -2766 -121620 -2366 -121580
rect -2047 -117450 -1647 -117410
rect -2047 -121580 -2007 -117450
rect -1687 -121580 -1647 -117450
rect -2047 -121620 -1647 -121580
rect -1328 -117450 -928 -117410
rect -1328 -121580 -1288 -117450
rect -968 -121580 -928 -117450
rect -1328 -121620 -928 -121580
rect -609 -117450 -209 -117410
rect -609 -121580 -569 -117450
rect -249 -121580 -209 -117450
rect -609 -121620 -209 -121580
rect 110 -117450 510 -117410
rect 110 -121580 150 -117450
rect 470 -121580 510 -117450
rect 110 -121620 510 -121580
rect 829 -117450 1229 -117410
rect 829 -121580 869 -117450
rect 1189 -121580 1229 -117450
rect 829 -121620 1229 -121580
rect 1548 -117450 1948 -117410
rect 1548 -121580 1588 -117450
rect 1908 -121580 1948 -117450
rect 1548 -121620 1948 -121580
rect 2267 -117450 2667 -117410
rect 2267 -121580 2307 -117450
rect 2627 -121580 2667 -117450
rect 2267 -121620 2667 -121580
rect -2766 -121960 -2366 -121920
rect -2766 -126090 -2726 -121960
rect -2406 -126090 -2366 -121960
rect -2766 -126130 -2366 -126090
rect -2047 -121960 -1647 -121920
rect -2047 -126090 -2007 -121960
rect -1687 -126090 -1647 -121960
rect -2047 -126130 -1647 -126090
rect -1328 -121960 -928 -121920
rect -1328 -126090 -1288 -121960
rect -968 -126090 -928 -121960
rect -1328 -126130 -928 -126090
rect -609 -121960 -209 -121920
rect -609 -126090 -569 -121960
rect -249 -126090 -209 -121960
rect -609 -126130 -209 -126090
rect 110 -121960 510 -121920
rect 110 -126090 150 -121960
rect 470 -126090 510 -121960
rect 110 -126130 510 -126090
rect 829 -121960 1229 -121920
rect 829 -126090 869 -121960
rect 1189 -126090 1229 -121960
rect 829 -126130 1229 -126090
rect 1548 -121960 1948 -121920
rect 1548 -126090 1588 -121960
rect 1908 -126090 1948 -121960
rect 1548 -126130 1948 -126090
rect 2267 -121960 2667 -121920
rect 2267 -126090 2307 -121960
rect 2627 -126090 2667 -121960
rect 2267 -126130 2667 -126090
rect -2766 -126470 -2366 -126430
rect -2766 -130600 -2726 -126470
rect -2406 -130600 -2366 -126470
rect -2766 -130640 -2366 -130600
rect -2047 -126470 -1647 -126430
rect -2047 -130600 -2007 -126470
rect -1687 -130600 -1647 -126470
rect -2047 -130640 -1647 -130600
rect -1328 -126470 -928 -126430
rect -1328 -130600 -1288 -126470
rect -968 -130600 -928 -126470
rect -1328 -130640 -928 -130600
rect -609 -126470 -209 -126430
rect -609 -130600 -569 -126470
rect -249 -130600 -209 -126470
rect -609 -130640 -209 -130600
rect 110 -126470 510 -126430
rect 110 -130600 150 -126470
rect 470 -130600 510 -126470
rect 110 -130640 510 -130600
rect 829 -126470 1229 -126430
rect 829 -130600 869 -126470
rect 1189 -130600 1229 -126470
rect 829 -130640 1229 -130600
rect 1548 -126470 1948 -126430
rect 1548 -130600 1588 -126470
rect 1908 -130600 1948 -126470
rect 1548 -130640 1948 -130600
rect 2267 -126470 2667 -126430
rect 2267 -130600 2307 -126470
rect 2627 -130600 2667 -126470
rect 2267 -130640 2667 -130600
rect -2766 -130980 -2366 -130940
rect -2766 -135110 -2726 -130980
rect -2406 -135110 -2366 -130980
rect -2766 -135150 -2366 -135110
rect -2047 -130980 -1647 -130940
rect -2047 -135110 -2007 -130980
rect -1687 -135110 -1647 -130980
rect -2047 -135150 -1647 -135110
rect -1328 -130980 -928 -130940
rect -1328 -135110 -1288 -130980
rect -968 -135110 -928 -130980
rect -1328 -135150 -928 -135110
rect -609 -130980 -209 -130940
rect -609 -135110 -569 -130980
rect -249 -135110 -209 -130980
rect -609 -135150 -209 -135110
rect 110 -130980 510 -130940
rect 110 -135110 150 -130980
rect 470 -135110 510 -130980
rect 110 -135150 510 -135110
rect 829 -130980 1229 -130940
rect 829 -135110 869 -130980
rect 1189 -135110 1229 -130980
rect 829 -135150 1229 -135110
rect 1548 -130980 1948 -130940
rect 1548 -135110 1588 -130980
rect 1908 -135110 1948 -130980
rect 1548 -135150 1948 -135110
rect 2267 -130980 2667 -130940
rect 2267 -135110 2307 -130980
rect 2627 -135110 2667 -130980
rect 2267 -135150 2667 -135110
rect -2766 -135490 -2366 -135450
rect -2766 -139620 -2726 -135490
rect -2406 -139620 -2366 -135490
rect -2766 -139660 -2366 -139620
rect -2047 -135490 -1647 -135450
rect -2047 -139620 -2007 -135490
rect -1687 -139620 -1647 -135490
rect -2047 -139660 -1647 -139620
rect -1328 -135490 -928 -135450
rect -1328 -139620 -1288 -135490
rect -968 -139620 -928 -135490
rect -1328 -139660 -928 -139620
rect -609 -135490 -209 -135450
rect -609 -139620 -569 -135490
rect -249 -139620 -209 -135490
rect -609 -139660 -209 -139620
rect 110 -135490 510 -135450
rect 110 -139620 150 -135490
rect 470 -139620 510 -135490
rect 110 -139660 510 -139620
rect 829 -135490 1229 -135450
rect 829 -139620 869 -135490
rect 1189 -139620 1229 -135490
rect 829 -139660 1229 -139620
rect 1548 -135490 1948 -135450
rect 1548 -139620 1588 -135490
rect 1908 -139620 1948 -135490
rect 1548 -139660 1948 -139620
rect 2267 -135490 2667 -135450
rect 2267 -139620 2307 -135490
rect 2627 -139620 2667 -135490
rect 2267 -139660 2667 -139620
rect -2766 -140000 -2366 -139960
rect -2766 -144130 -2726 -140000
rect -2406 -144130 -2366 -140000
rect -2766 -144170 -2366 -144130
rect -2047 -140000 -1647 -139960
rect -2047 -144130 -2007 -140000
rect -1687 -144130 -1647 -140000
rect -2047 -144170 -1647 -144130
rect -1328 -140000 -928 -139960
rect -1328 -144130 -1288 -140000
rect -968 -144130 -928 -140000
rect -1328 -144170 -928 -144130
rect -609 -140000 -209 -139960
rect -609 -144130 -569 -140000
rect -249 -144130 -209 -140000
rect -609 -144170 -209 -144130
rect 110 -140000 510 -139960
rect 110 -144130 150 -140000
rect 470 -144130 510 -140000
rect 110 -144170 510 -144130
rect 829 -140000 1229 -139960
rect 829 -144130 869 -140000
rect 1189 -144130 1229 -140000
rect 829 -144170 1229 -144130
rect 1548 -140000 1948 -139960
rect 1548 -144130 1588 -140000
rect 1908 -144130 1948 -140000
rect 1548 -144170 1948 -144130
rect 2267 -140000 2667 -139960
rect 2267 -144130 2307 -140000
rect 2627 -144130 2667 -140000
rect 2267 -144170 2667 -144130
<< mimcapcontact >>
rect -2726 140000 -2406 144130
rect -2007 140000 -1687 144130
rect -1288 140000 -968 144130
rect -569 140000 -249 144130
rect 150 140000 470 144130
rect 869 140000 1189 144130
rect 1588 140000 1908 144130
rect 2307 140000 2627 144130
rect -2726 135490 -2406 139620
rect -2007 135490 -1687 139620
rect -1288 135490 -968 139620
rect -569 135490 -249 139620
rect 150 135490 470 139620
rect 869 135490 1189 139620
rect 1588 135490 1908 139620
rect 2307 135490 2627 139620
rect -2726 130980 -2406 135110
rect -2007 130980 -1687 135110
rect -1288 130980 -968 135110
rect -569 130980 -249 135110
rect 150 130980 470 135110
rect 869 130980 1189 135110
rect 1588 130980 1908 135110
rect 2307 130980 2627 135110
rect -2726 126470 -2406 130600
rect -2007 126470 -1687 130600
rect -1288 126470 -968 130600
rect -569 126470 -249 130600
rect 150 126470 470 130600
rect 869 126470 1189 130600
rect 1588 126470 1908 130600
rect 2307 126470 2627 130600
rect -2726 121960 -2406 126090
rect -2007 121960 -1687 126090
rect -1288 121960 -968 126090
rect -569 121960 -249 126090
rect 150 121960 470 126090
rect 869 121960 1189 126090
rect 1588 121960 1908 126090
rect 2307 121960 2627 126090
rect -2726 117450 -2406 121580
rect -2007 117450 -1687 121580
rect -1288 117450 -968 121580
rect -569 117450 -249 121580
rect 150 117450 470 121580
rect 869 117450 1189 121580
rect 1588 117450 1908 121580
rect 2307 117450 2627 121580
rect -2726 112940 -2406 117070
rect -2007 112940 -1687 117070
rect -1288 112940 -968 117070
rect -569 112940 -249 117070
rect 150 112940 470 117070
rect 869 112940 1189 117070
rect 1588 112940 1908 117070
rect 2307 112940 2627 117070
rect -2726 108430 -2406 112560
rect -2007 108430 -1687 112560
rect -1288 108430 -968 112560
rect -569 108430 -249 112560
rect 150 108430 470 112560
rect 869 108430 1189 112560
rect 1588 108430 1908 112560
rect 2307 108430 2627 112560
rect -2726 103920 -2406 108050
rect -2007 103920 -1687 108050
rect -1288 103920 -968 108050
rect -569 103920 -249 108050
rect 150 103920 470 108050
rect 869 103920 1189 108050
rect 1588 103920 1908 108050
rect 2307 103920 2627 108050
rect -2726 99410 -2406 103540
rect -2007 99410 -1687 103540
rect -1288 99410 -968 103540
rect -569 99410 -249 103540
rect 150 99410 470 103540
rect 869 99410 1189 103540
rect 1588 99410 1908 103540
rect 2307 99410 2627 103540
rect -2726 94900 -2406 99030
rect -2007 94900 -1687 99030
rect -1288 94900 -968 99030
rect -569 94900 -249 99030
rect 150 94900 470 99030
rect 869 94900 1189 99030
rect 1588 94900 1908 99030
rect 2307 94900 2627 99030
rect -2726 90390 -2406 94520
rect -2007 90390 -1687 94520
rect -1288 90390 -968 94520
rect -569 90390 -249 94520
rect 150 90390 470 94520
rect 869 90390 1189 94520
rect 1588 90390 1908 94520
rect 2307 90390 2627 94520
rect -2726 85880 -2406 90010
rect -2007 85880 -1687 90010
rect -1288 85880 -968 90010
rect -569 85880 -249 90010
rect 150 85880 470 90010
rect 869 85880 1189 90010
rect 1588 85880 1908 90010
rect 2307 85880 2627 90010
rect -2726 81370 -2406 85500
rect -2007 81370 -1687 85500
rect -1288 81370 -968 85500
rect -569 81370 -249 85500
rect 150 81370 470 85500
rect 869 81370 1189 85500
rect 1588 81370 1908 85500
rect 2307 81370 2627 85500
rect -2726 76860 -2406 80990
rect -2007 76860 -1687 80990
rect -1288 76860 -968 80990
rect -569 76860 -249 80990
rect 150 76860 470 80990
rect 869 76860 1189 80990
rect 1588 76860 1908 80990
rect 2307 76860 2627 80990
rect -2726 72350 -2406 76480
rect -2007 72350 -1687 76480
rect -1288 72350 -968 76480
rect -569 72350 -249 76480
rect 150 72350 470 76480
rect 869 72350 1189 76480
rect 1588 72350 1908 76480
rect 2307 72350 2627 76480
rect -2726 67840 -2406 71970
rect -2007 67840 -1687 71970
rect -1288 67840 -968 71970
rect -569 67840 -249 71970
rect 150 67840 470 71970
rect 869 67840 1189 71970
rect 1588 67840 1908 71970
rect 2307 67840 2627 71970
rect -2726 63330 -2406 67460
rect -2007 63330 -1687 67460
rect -1288 63330 -968 67460
rect -569 63330 -249 67460
rect 150 63330 470 67460
rect 869 63330 1189 67460
rect 1588 63330 1908 67460
rect 2307 63330 2627 67460
rect -2726 58820 -2406 62950
rect -2007 58820 -1687 62950
rect -1288 58820 -968 62950
rect -569 58820 -249 62950
rect 150 58820 470 62950
rect 869 58820 1189 62950
rect 1588 58820 1908 62950
rect 2307 58820 2627 62950
rect -2726 54310 -2406 58440
rect -2007 54310 -1687 58440
rect -1288 54310 -968 58440
rect -569 54310 -249 58440
rect 150 54310 470 58440
rect 869 54310 1189 58440
rect 1588 54310 1908 58440
rect 2307 54310 2627 58440
rect -2726 49800 -2406 53930
rect -2007 49800 -1687 53930
rect -1288 49800 -968 53930
rect -569 49800 -249 53930
rect 150 49800 470 53930
rect 869 49800 1189 53930
rect 1588 49800 1908 53930
rect 2307 49800 2627 53930
rect -2726 45290 -2406 49420
rect -2007 45290 -1687 49420
rect -1288 45290 -968 49420
rect -569 45290 -249 49420
rect 150 45290 470 49420
rect 869 45290 1189 49420
rect 1588 45290 1908 49420
rect 2307 45290 2627 49420
rect -2726 40780 -2406 44910
rect -2007 40780 -1687 44910
rect -1288 40780 -968 44910
rect -569 40780 -249 44910
rect 150 40780 470 44910
rect 869 40780 1189 44910
rect 1588 40780 1908 44910
rect 2307 40780 2627 44910
rect -2726 36270 -2406 40400
rect -2007 36270 -1687 40400
rect -1288 36270 -968 40400
rect -569 36270 -249 40400
rect 150 36270 470 40400
rect 869 36270 1189 40400
rect 1588 36270 1908 40400
rect 2307 36270 2627 40400
rect -2726 31760 -2406 35890
rect -2007 31760 -1687 35890
rect -1288 31760 -968 35890
rect -569 31760 -249 35890
rect 150 31760 470 35890
rect 869 31760 1189 35890
rect 1588 31760 1908 35890
rect 2307 31760 2627 35890
rect -2726 27250 -2406 31380
rect -2007 27250 -1687 31380
rect -1288 27250 -968 31380
rect -569 27250 -249 31380
rect 150 27250 470 31380
rect 869 27250 1189 31380
rect 1588 27250 1908 31380
rect 2307 27250 2627 31380
rect -2726 22740 -2406 26870
rect -2007 22740 -1687 26870
rect -1288 22740 -968 26870
rect -569 22740 -249 26870
rect 150 22740 470 26870
rect 869 22740 1189 26870
rect 1588 22740 1908 26870
rect 2307 22740 2627 26870
rect -2726 18230 -2406 22360
rect -2007 18230 -1687 22360
rect -1288 18230 -968 22360
rect -569 18230 -249 22360
rect 150 18230 470 22360
rect 869 18230 1189 22360
rect 1588 18230 1908 22360
rect 2307 18230 2627 22360
rect -2726 13720 -2406 17850
rect -2007 13720 -1687 17850
rect -1288 13720 -968 17850
rect -569 13720 -249 17850
rect 150 13720 470 17850
rect 869 13720 1189 17850
rect 1588 13720 1908 17850
rect 2307 13720 2627 17850
rect -2726 9210 -2406 13340
rect -2007 9210 -1687 13340
rect -1288 9210 -968 13340
rect -569 9210 -249 13340
rect 150 9210 470 13340
rect 869 9210 1189 13340
rect 1588 9210 1908 13340
rect 2307 9210 2627 13340
rect -2726 4700 -2406 8830
rect -2007 4700 -1687 8830
rect -1288 4700 -968 8830
rect -569 4700 -249 8830
rect 150 4700 470 8830
rect 869 4700 1189 8830
rect 1588 4700 1908 8830
rect 2307 4700 2627 8830
rect -2726 190 -2406 4320
rect -2007 190 -1687 4320
rect -1288 190 -968 4320
rect -569 190 -249 4320
rect 150 190 470 4320
rect 869 190 1189 4320
rect 1588 190 1908 4320
rect 2307 190 2627 4320
rect -2726 -4320 -2406 -190
rect -2007 -4320 -1687 -190
rect -1288 -4320 -968 -190
rect -569 -4320 -249 -190
rect 150 -4320 470 -190
rect 869 -4320 1189 -190
rect 1588 -4320 1908 -190
rect 2307 -4320 2627 -190
rect -2726 -8830 -2406 -4700
rect -2007 -8830 -1687 -4700
rect -1288 -8830 -968 -4700
rect -569 -8830 -249 -4700
rect 150 -8830 470 -4700
rect 869 -8830 1189 -4700
rect 1588 -8830 1908 -4700
rect 2307 -8830 2627 -4700
rect -2726 -13340 -2406 -9210
rect -2007 -13340 -1687 -9210
rect -1288 -13340 -968 -9210
rect -569 -13340 -249 -9210
rect 150 -13340 470 -9210
rect 869 -13340 1189 -9210
rect 1588 -13340 1908 -9210
rect 2307 -13340 2627 -9210
rect -2726 -17850 -2406 -13720
rect -2007 -17850 -1687 -13720
rect -1288 -17850 -968 -13720
rect -569 -17850 -249 -13720
rect 150 -17850 470 -13720
rect 869 -17850 1189 -13720
rect 1588 -17850 1908 -13720
rect 2307 -17850 2627 -13720
rect -2726 -22360 -2406 -18230
rect -2007 -22360 -1687 -18230
rect -1288 -22360 -968 -18230
rect -569 -22360 -249 -18230
rect 150 -22360 470 -18230
rect 869 -22360 1189 -18230
rect 1588 -22360 1908 -18230
rect 2307 -22360 2627 -18230
rect -2726 -26870 -2406 -22740
rect -2007 -26870 -1687 -22740
rect -1288 -26870 -968 -22740
rect -569 -26870 -249 -22740
rect 150 -26870 470 -22740
rect 869 -26870 1189 -22740
rect 1588 -26870 1908 -22740
rect 2307 -26870 2627 -22740
rect -2726 -31380 -2406 -27250
rect -2007 -31380 -1687 -27250
rect -1288 -31380 -968 -27250
rect -569 -31380 -249 -27250
rect 150 -31380 470 -27250
rect 869 -31380 1189 -27250
rect 1588 -31380 1908 -27250
rect 2307 -31380 2627 -27250
rect -2726 -35890 -2406 -31760
rect -2007 -35890 -1687 -31760
rect -1288 -35890 -968 -31760
rect -569 -35890 -249 -31760
rect 150 -35890 470 -31760
rect 869 -35890 1189 -31760
rect 1588 -35890 1908 -31760
rect 2307 -35890 2627 -31760
rect -2726 -40400 -2406 -36270
rect -2007 -40400 -1687 -36270
rect -1288 -40400 -968 -36270
rect -569 -40400 -249 -36270
rect 150 -40400 470 -36270
rect 869 -40400 1189 -36270
rect 1588 -40400 1908 -36270
rect 2307 -40400 2627 -36270
rect -2726 -44910 -2406 -40780
rect -2007 -44910 -1687 -40780
rect -1288 -44910 -968 -40780
rect -569 -44910 -249 -40780
rect 150 -44910 470 -40780
rect 869 -44910 1189 -40780
rect 1588 -44910 1908 -40780
rect 2307 -44910 2627 -40780
rect -2726 -49420 -2406 -45290
rect -2007 -49420 -1687 -45290
rect -1288 -49420 -968 -45290
rect -569 -49420 -249 -45290
rect 150 -49420 470 -45290
rect 869 -49420 1189 -45290
rect 1588 -49420 1908 -45290
rect 2307 -49420 2627 -45290
rect -2726 -53930 -2406 -49800
rect -2007 -53930 -1687 -49800
rect -1288 -53930 -968 -49800
rect -569 -53930 -249 -49800
rect 150 -53930 470 -49800
rect 869 -53930 1189 -49800
rect 1588 -53930 1908 -49800
rect 2307 -53930 2627 -49800
rect -2726 -58440 -2406 -54310
rect -2007 -58440 -1687 -54310
rect -1288 -58440 -968 -54310
rect -569 -58440 -249 -54310
rect 150 -58440 470 -54310
rect 869 -58440 1189 -54310
rect 1588 -58440 1908 -54310
rect 2307 -58440 2627 -54310
rect -2726 -62950 -2406 -58820
rect -2007 -62950 -1687 -58820
rect -1288 -62950 -968 -58820
rect -569 -62950 -249 -58820
rect 150 -62950 470 -58820
rect 869 -62950 1189 -58820
rect 1588 -62950 1908 -58820
rect 2307 -62950 2627 -58820
rect -2726 -67460 -2406 -63330
rect -2007 -67460 -1687 -63330
rect -1288 -67460 -968 -63330
rect -569 -67460 -249 -63330
rect 150 -67460 470 -63330
rect 869 -67460 1189 -63330
rect 1588 -67460 1908 -63330
rect 2307 -67460 2627 -63330
rect -2726 -71970 -2406 -67840
rect -2007 -71970 -1687 -67840
rect -1288 -71970 -968 -67840
rect -569 -71970 -249 -67840
rect 150 -71970 470 -67840
rect 869 -71970 1189 -67840
rect 1588 -71970 1908 -67840
rect 2307 -71970 2627 -67840
rect -2726 -76480 -2406 -72350
rect -2007 -76480 -1687 -72350
rect -1288 -76480 -968 -72350
rect -569 -76480 -249 -72350
rect 150 -76480 470 -72350
rect 869 -76480 1189 -72350
rect 1588 -76480 1908 -72350
rect 2307 -76480 2627 -72350
rect -2726 -80990 -2406 -76860
rect -2007 -80990 -1687 -76860
rect -1288 -80990 -968 -76860
rect -569 -80990 -249 -76860
rect 150 -80990 470 -76860
rect 869 -80990 1189 -76860
rect 1588 -80990 1908 -76860
rect 2307 -80990 2627 -76860
rect -2726 -85500 -2406 -81370
rect -2007 -85500 -1687 -81370
rect -1288 -85500 -968 -81370
rect -569 -85500 -249 -81370
rect 150 -85500 470 -81370
rect 869 -85500 1189 -81370
rect 1588 -85500 1908 -81370
rect 2307 -85500 2627 -81370
rect -2726 -90010 -2406 -85880
rect -2007 -90010 -1687 -85880
rect -1288 -90010 -968 -85880
rect -569 -90010 -249 -85880
rect 150 -90010 470 -85880
rect 869 -90010 1189 -85880
rect 1588 -90010 1908 -85880
rect 2307 -90010 2627 -85880
rect -2726 -94520 -2406 -90390
rect -2007 -94520 -1687 -90390
rect -1288 -94520 -968 -90390
rect -569 -94520 -249 -90390
rect 150 -94520 470 -90390
rect 869 -94520 1189 -90390
rect 1588 -94520 1908 -90390
rect 2307 -94520 2627 -90390
rect -2726 -99030 -2406 -94900
rect -2007 -99030 -1687 -94900
rect -1288 -99030 -968 -94900
rect -569 -99030 -249 -94900
rect 150 -99030 470 -94900
rect 869 -99030 1189 -94900
rect 1588 -99030 1908 -94900
rect 2307 -99030 2627 -94900
rect -2726 -103540 -2406 -99410
rect -2007 -103540 -1687 -99410
rect -1288 -103540 -968 -99410
rect -569 -103540 -249 -99410
rect 150 -103540 470 -99410
rect 869 -103540 1189 -99410
rect 1588 -103540 1908 -99410
rect 2307 -103540 2627 -99410
rect -2726 -108050 -2406 -103920
rect -2007 -108050 -1687 -103920
rect -1288 -108050 -968 -103920
rect -569 -108050 -249 -103920
rect 150 -108050 470 -103920
rect 869 -108050 1189 -103920
rect 1588 -108050 1908 -103920
rect 2307 -108050 2627 -103920
rect -2726 -112560 -2406 -108430
rect -2007 -112560 -1687 -108430
rect -1288 -112560 -968 -108430
rect -569 -112560 -249 -108430
rect 150 -112560 470 -108430
rect 869 -112560 1189 -108430
rect 1588 -112560 1908 -108430
rect 2307 -112560 2627 -108430
rect -2726 -117070 -2406 -112940
rect -2007 -117070 -1687 -112940
rect -1288 -117070 -968 -112940
rect -569 -117070 -249 -112940
rect 150 -117070 470 -112940
rect 869 -117070 1189 -112940
rect 1588 -117070 1908 -112940
rect 2307 -117070 2627 -112940
rect -2726 -121580 -2406 -117450
rect -2007 -121580 -1687 -117450
rect -1288 -121580 -968 -117450
rect -569 -121580 -249 -117450
rect 150 -121580 470 -117450
rect 869 -121580 1189 -117450
rect 1588 -121580 1908 -117450
rect 2307 -121580 2627 -117450
rect -2726 -126090 -2406 -121960
rect -2007 -126090 -1687 -121960
rect -1288 -126090 -968 -121960
rect -569 -126090 -249 -121960
rect 150 -126090 470 -121960
rect 869 -126090 1189 -121960
rect 1588 -126090 1908 -121960
rect 2307 -126090 2627 -121960
rect -2726 -130600 -2406 -126470
rect -2007 -130600 -1687 -126470
rect -1288 -130600 -968 -126470
rect -569 -130600 -249 -126470
rect 150 -130600 470 -126470
rect 869 -130600 1189 -126470
rect 1588 -130600 1908 -126470
rect 2307 -130600 2627 -126470
rect -2726 -135110 -2406 -130980
rect -2007 -135110 -1687 -130980
rect -1288 -135110 -968 -130980
rect -569 -135110 -249 -130980
rect 150 -135110 470 -130980
rect 869 -135110 1189 -130980
rect 1588 -135110 1908 -130980
rect 2307 -135110 2627 -130980
rect -2726 -139620 -2406 -135490
rect -2007 -139620 -1687 -135490
rect -1288 -139620 -968 -135490
rect -569 -139620 -249 -135490
rect 150 -139620 470 -135490
rect 869 -139620 1189 -135490
rect 1588 -139620 1908 -135490
rect 2307 -139620 2627 -135490
rect -2726 -144130 -2406 -140000
rect -2007 -144130 -1687 -140000
rect -1288 -144130 -968 -140000
rect -569 -144130 -249 -140000
rect 150 -144130 470 -140000
rect 869 -144130 1189 -140000
rect 1588 -144130 1908 -140000
rect 2307 -144130 2627 -140000
<< metal4 >>
rect -2618 144131 -2514 144320
rect -2298 144258 -2194 144320
rect -2298 144242 -2171 144258
rect -2727 144130 -2405 144131
rect -2727 140000 -2726 144130
rect -2406 140000 -2405 144130
rect -2727 139999 -2405 140000
rect -2618 139621 -2514 139999
rect -2298 139888 -2251 144242
rect -2187 139888 -2171 144242
rect -1899 144131 -1795 144320
rect -1579 144258 -1475 144320
rect -1579 144242 -1452 144258
rect -2008 144130 -1686 144131
rect -2008 140000 -2007 144130
rect -1687 140000 -1686 144130
rect -2008 139999 -1686 140000
rect -2298 139872 -2171 139888
rect -2298 139748 -2194 139872
rect -2298 139732 -2171 139748
rect -2727 139620 -2405 139621
rect -2727 135490 -2726 139620
rect -2406 135490 -2405 139620
rect -2727 135489 -2405 135490
rect -2618 135111 -2514 135489
rect -2298 135378 -2251 139732
rect -2187 135378 -2171 139732
rect -1899 139621 -1795 139999
rect -1579 139888 -1532 144242
rect -1468 139888 -1452 144242
rect -1180 144131 -1076 144320
rect -860 144258 -756 144320
rect -860 144242 -733 144258
rect -1289 144130 -967 144131
rect -1289 140000 -1288 144130
rect -968 140000 -967 144130
rect -1289 139999 -967 140000
rect -1579 139872 -1452 139888
rect -1579 139748 -1475 139872
rect -1579 139732 -1452 139748
rect -2008 139620 -1686 139621
rect -2008 135490 -2007 139620
rect -1687 135490 -1686 139620
rect -2008 135489 -1686 135490
rect -2298 135362 -2171 135378
rect -2298 135238 -2194 135362
rect -2298 135222 -2171 135238
rect -2727 135110 -2405 135111
rect -2727 130980 -2726 135110
rect -2406 130980 -2405 135110
rect -2727 130979 -2405 130980
rect -2618 130601 -2514 130979
rect -2298 130868 -2251 135222
rect -2187 130868 -2171 135222
rect -1899 135111 -1795 135489
rect -1579 135378 -1532 139732
rect -1468 135378 -1452 139732
rect -1180 139621 -1076 139999
rect -860 139888 -813 144242
rect -749 139888 -733 144242
rect -461 144131 -357 144320
rect -141 144258 -37 144320
rect -141 144242 -14 144258
rect -570 144130 -248 144131
rect -570 140000 -569 144130
rect -249 140000 -248 144130
rect -570 139999 -248 140000
rect -860 139872 -733 139888
rect -860 139748 -756 139872
rect -860 139732 -733 139748
rect -1289 139620 -967 139621
rect -1289 135490 -1288 139620
rect -968 135490 -967 139620
rect -1289 135489 -967 135490
rect -1579 135362 -1452 135378
rect -1579 135238 -1475 135362
rect -1579 135222 -1452 135238
rect -2008 135110 -1686 135111
rect -2008 130980 -2007 135110
rect -1687 130980 -1686 135110
rect -2008 130979 -1686 130980
rect -2298 130852 -2171 130868
rect -2298 130728 -2194 130852
rect -2298 130712 -2171 130728
rect -2727 130600 -2405 130601
rect -2727 126470 -2726 130600
rect -2406 126470 -2405 130600
rect -2727 126469 -2405 126470
rect -2618 126091 -2514 126469
rect -2298 126358 -2251 130712
rect -2187 126358 -2171 130712
rect -1899 130601 -1795 130979
rect -1579 130868 -1532 135222
rect -1468 130868 -1452 135222
rect -1180 135111 -1076 135489
rect -860 135378 -813 139732
rect -749 135378 -733 139732
rect -461 139621 -357 139999
rect -141 139888 -94 144242
rect -30 139888 -14 144242
rect 258 144131 362 144320
rect 578 144258 682 144320
rect 578 144242 705 144258
rect 149 144130 471 144131
rect 149 140000 150 144130
rect 470 140000 471 144130
rect 149 139999 471 140000
rect -141 139872 -14 139888
rect -141 139748 -37 139872
rect -141 139732 -14 139748
rect -570 139620 -248 139621
rect -570 135490 -569 139620
rect -249 135490 -248 139620
rect -570 135489 -248 135490
rect -860 135362 -733 135378
rect -860 135238 -756 135362
rect -860 135222 -733 135238
rect -1289 135110 -967 135111
rect -1289 130980 -1288 135110
rect -968 130980 -967 135110
rect -1289 130979 -967 130980
rect -1579 130852 -1452 130868
rect -1579 130728 -1475 130852
rect -1579 130712 -1452 130728
rect -2008 130600 -1686 130601
rect -2008 126470 -2007 130600
rect -1687 126470 -1686 130600
rect -2008 126469 -1686 126470
rect -2298 126342 -2171 126358
rect -2298 126218 -2194 126342
rect -2298 126202 -2171 126218
rect -2727 126090 -2405 126091
rect -2727 121960 -2726 126090
rect -2406 121960 -2405 126090
rect -2727 121959 -2405 121960
rect -2618 121581 -2514 121959
rect -2298 121848 -2251 126202
rect -2187 121848 -2171 126202
rect -1899 126091 -1795 126469
rect -1579 126358 -1532 130712
rect -1468 126358 -1452 130712
rect -1180 130601 -1076 130979
rect -860 130868 -813 135222
rect -749 130868 -733 135222
rect -461 135111 -357 135489
rect -141 135378 -94 139732
rect -30 135378 -14 139732
rect 258 139621 362 139999
rect 578 139888 625 144242
rect 689 139888 705 144242
rect 977 144131 1081 144320
rect 1297 144258 1401 144320
rect 1297 144242 1424 144258
rect 868 144130 1190 144131
rect 868 140000 869 144130
rect 1189 140000 1190 144130
rect 868 139999 1190 140000
rect 578 139872 705 139888
rect 578 139748 682 139872
rect 578 139732 705 139748
rect 149 139620 471 139621
rect 149 135490 150 139620
rect 470 135490 471 139620
rect 149 135489 471 135490
rect -141 135362 -14 135378
rect -141 135238 -37 135362
rect -141 135222 -14 135238
rect -570 135110 -248 135111
rect -570 130980 -569 135110
rect -249 130980 -248 135110
rect -570 130979 -248 130980
rect -860 130852 -733 130868
rect -860 130728 -756 130852
rect -860 130712 -733 130728
rect -1289 130600 -967 130601
rect -1289 126470 -1288 130600
rect -968 126470 -967 130600
rect -1289 126469 -967 126470
rect -1579 126342 -1452 126358
rect -1579 126218 -1475 126342
rect -1579 126202 -1452 126218
rect -2008 126090 -1686 126091
rect -2008 121960 -2007 126090
rect -1687 121960 -1686 126090
rect -2008 121959 -1686 121960
rect -2298 121832 -2171 121848
rect -2298 121708 -2194 121832
rect -2298 121692 -2171 121708
rect -2727 121580 -2405 121581
rect -2727 117450 -2726 121580
rect -2406 117450 -2405 121580
rect -2727 117449 -2405 117450
rect -2618 117071 -2514 117449
rect -2298 117338 -2251 121692
rect -2187 117338 -2171 121692
rect -1899 121581 -1795 121959
rect -1579 121848 -1532 126202
rect -1468 121848 -1452 126202
rect -1180 126091 -1076 126469
rect -860 126358 -813 130712
rect -749 126358 -733 130712
rect -461 130601 -357 130979
rect -141 130868 -94 135222
rect -30 130868 -14 135222
rect 258 135111 362 135489
rect 578 135378 625 139732
rect 689 135378 705 139732
rect 977 139621 1081 139999
rect 1297 139888 1344 144242
rect 1408 139888 1424 144242
rect 1696 144131 1800 144320
rect 2016 144258 2120 144320
rect 2016 144242 2143 144258
rect 1587 144130 1909 144131
rect 1587 140000 1588 144130
rect 1908 140000 1909 144130
rect 1587 139999 1909 140000
rect 1297 139872 1424 139888
rect 1297 139748 1401 139872
rect 1297 139732 1424 139748
rect 868 139620 1190 139621
rect 868 135490 869 139620
rect 1189 135490 1190 139620
rect 868 135489 1190 135490
rect 578 135362 705 135378
rect 578 135238 682 135362
rect 578 135222 705 135238
rect 149 135110 471 135111
rect 149 130980 150 135110
rect 470 130980 471 135110
rect 149 130979 471 130980
rect -141 130852 -14 130868
rect -141 130728 -37 130852
rect -141 130712 -14 130728
rect -570 130600 -248 130601
rect -570 126470 -569 130600
rect -249 126470 -248 130600
rect -570 126469 -248 126470
rect -860 126342 -733 126358
rect -860 126218 -756 126342
rect -860 126202 -733 126218
rect -1289 126090 -967 126091
rect -1289 121960 -1288 126090
rect -968 121960 -967 126090
rect -1289 121959 -967 121960
rect -1579 121832 -1452 121848
rect -1579 121708 -1475 121832
rect -1579 121692 -1452 121708
rect -2008 121580 -1686 121581
rect -2008 117450 -2007 121580
rect -1687 117450 -1686 121580
rect -2008 117449 -1686 117450
rect -2298 117322 -2171 117338
rect -2298 117198 -2194 117322
rect -2298 117182 -2171 117198
rect -2727 117070 -2405 117071
rect -2727 112940 -2726 117070
rect -2406 112940 -2405 117070
rect -2727 112939 -2405 112940
rect -2618 112561 -2514 112939
rect -2298 112828 -2251 117182
rect -2187 112828 -2171 117182
rect -1899 117071 -1795 117449
rect -1579 117338 -1532 121692
rect -1468 117338 -1452 121692
rect -1180 121581 -1076 121959
rect -860 121848 -813 126202
rect -749 121848 -733 126202
rect -461 126091 -357 126469
rect -141 126358 -94 130712
rect -30 126358 -14 130712
rect 258 130601 362 130979
rect 578 130868 625 135222
rect 689 130868 705 135222
rect 977 135111 1081 135489
rect 1297 135378 1344 139732
rect 1408 135378 1424 139732
rect 1696 139621 1800 139999
rect 2016 139888 2063 144242
rect 2127 139888 2143 144242
rect 2415 144131 2519 144320
rect 2735 144258 2839 144320
rect 2735 144242 2862 144258
rect 2306 144130 2628 144131
rect 2306 140000 2307 144130
rect 2627 140000 2628 144130
rect 2306 139999 2628 140000
rect 2016 139872 2143 139888
rect 2016 139748 2120 139872
rect 2016 139732 2143 139748
rect 1587 139620 1909 139621
rect 1587 135490 1588 139620
rect 1908 135490 1909 139620
rect 1587 135489 1909 135490
rect 1297 135362 1424 135378
rect 1297 135238 1401 135362
rect 1297 135222 1424 135238
rect 868 135110 1190 135111
rect 868 130980 869 135110
rect 1189 130980 1190 135110
rect 868 130979 1190 130980
rect 578 130852 705 130868
rect 578 130728 682 130852
rect 578 130712 705 130728
rect 149 130600 471 130601
rect 149 126470 150 130600
rect 470 126470 471 130600
rect 149 126469 471 126470
rect -141 126342 -14 126358
rect -141 126218 -37 126342
rect -141 126202 -14 126218
rect -570 126090 -248 126091
rect -570 121960 -569 126090
rect -249 121960 -248 126090
rect -570 121959 -248 121960
rect -860 121832 -733 121848
rect -860 121708 -756 121832
rect -860 121692 -733 121708
rect -1289 121580 -967 121581
rect -1289 117450 -1288 121580
rect -968 117450 -967 121580
rect -1289 117449 -967 117450
rect -1579 117322 -1452 117338
rect -1579 117198 -1475 117322
rect -1579 117182 -1452 117198
rect -2008 117070 -1686 117071
rect -2008 112940 -2007 117070
rect -1687 112940 -1686 117070
rect -2008 112939 -1686 112940
rect -2298 112812 -2171 112828
rect -2298 112688 -2194 112812
rect -2298 112672 -2171 112688
rect -2727 112560 -2405 112561
rect -2727 108430 -2726 112560
rect -2406 108430 -2405 112560
rect -2727 108429 -2405 108430
rect -2618 108051 -2514 108429
rect -2298 108318 -2251 112672
rect -2187 108318 -2171 112672
rect -1899 112561 -1795 112939
rect -1579 112828 -1532 117182
rect -1468 112828 -1452 117182
rect -1180 117071 -1076 117449
rect -860 117338 -813 121692
rect -749 117338 -733 121692
rect -461 121581 -357 121959
rect -141 121848 -94 126202
rect -30 121848 -14 126202
rect 258 126091 362 126469
rect 578 126358 625 130712
rect 689 126358 705 130712
rect 977 130601 1081 130979
rect 1297 130868 1344 135222
rect 1408 130868 1424 135222
rect 1696 135111 1800 135489
rect 2016 135378 2063 139732
rect 2127 135378 2143 139732
rect 2415 139621 2519 139999
rect 2735 139888 2782 144242
rect 2846 139888 2862 144242
rect 2735 139872 2862 139888
rect 2735 139748 2839 139872
rect 2735 139732 2862 139748
rect 2306 139620 2628 139621
rect 2306 135490 2307 139620
rect 2627 135490 2628 139620
rect 2306 135489 2628 135490
rect 2016 135362 2143 135378
rect 2016 135238 2120 135362
rect 2016 135222 2143 135238
rect 1587 135110 1909 135111
rect 1587 130980 1588 135110
rect 1908 130980 1909 135110
rect 1587 130979 1909 130980
rect 1297 130852 1424 130868
rect 1297 130728 1401 130852
rect 1297 130712 1424 130728
rect 868 130600 1190 130601
rect 868 126470 869 130600
rect 1189 126470 1190 130600
rect 868 126469 1190 126470
rect 578 126342 705 126358
rect 578 126218 682 126342
rect 578 126202 705 126218
rect 149 126090 471 126091
rect 149 121960 150 126090
rect 470 121960 471 126090
rect 149 121959 471 121960
rect -141 121832 -14 121848
rect -141 121708 -37 121832
rect -141 121692 -14 121708
rect -570 121580 -248 121581
rect -570 117450 -569 121580
rect -249 117450 -248 121580
rect -570 117449 -248 117450
rect -860 117322 -733 117338
rect -860 117198 -756 117322
rect -860 117182 -733 117198
rect -1289 117070 -967 117071
rect -1289 112940 -1288 117070
rect -968 112940 -967 117070
rect -1289 112939 -967 112940
rect -1579 112812 -1452 112828
rect -1579 112688 -1475 112812
rect -1579 112672 -1452 112688
rect -2008 112560 -1686 112561
rect -2008 108430 -2007 112560
rect -1687 108430 -1686 112560
rect -2008 108429 -1686 108430
rect -2298 108302 -2171 108318
rect -2298 108178 -2194 108302
rect -2298 108162 -2171 108178
rect -2727 108050 -2405 108051
rect -2727 103920 -2726 108050
rect -2406 103920 -2405 108050
rect -2727 103919 -2405 103920
rect -2618 103541 -2514 103919
rect -2298 103808 -2251 108162
rect -2187 103808 -2171 108162
rect -1899 108051 -1795 108429
rect -1579 108318 -1532 112672
rect -1468 108318 -1452 112672
rect -1180 112561 -1076 112939
rect -860 112828 -813 117182
rect -749 112828 -733 117182
rect -461 117071 -357 117449
rect -141 117338 -94 121692
rect -30 117338 -14 121692
rect 258 121581 362 121959
rect 578 121848 625 126202
rect 689 121848 705 126202
rect 977 126091 1081 126469
rect 1297 126358 1344 130712
rect 1408 126358 1424 130712
rect 1696 130601 1800 130979
rect 2016 130868 2063 135222
rect 2127 130868 2143 135222
rect 2415 135111 2519 135489
rect 2735 135378 2782 139732
rect 2846 135378 2862 139732
rect 2735 135362 2862 135378
rect 2735 135238 2839 135362
rect 2735 135222 2862 135238
rect 2306 135110 2628 135111
rect 2306 130980 2307 135110
rect 2627 130980 2628 135110
rect 2306 130979 2628 130980
rect 2016 130852 2143 130868
rect 2016 130728 2120 130852
rect 2016 130712 2143 130728
rect 1587 130600 1909 130601
rect 1587 126470 1588 130600
rect 1908 126470 1909 130600
rect 1587 126469 1909 126470
rect 1297 126342 1424 126358
rect 1297 126218 1401 126342
rect 1297 126202 1424 126218
rect 868 126090 1190 126091
rect 868 121960 869 126090
rect 1189 121960 1190 126090
rect 868 121959 1190 121960
rect 578 121832 705 121848
rect 578 121708 682 121832
rect 578 121692 705 121708
rect 149 121580 471 121581
rect 149 117450 150 121580
rect 470 117450 471 121580
rect 149 117449 471 117450
rect -141 117322 -14 117338
rect -141 117198 -37 117322
rect -141 117182 -14 117198
rect -570 117070 -248 117071
rect -570 112940 -569 117070
rect -249 112940 -248 117070
rect -570 112939 -248 112940
rect -860 112812 -733 112828
rect -860 112688 -756 112812
rect -860 112672 -733 112688
rect -1289 112560 -967 112561
rect -1289 108430 -1288 112560
rect -968 108430 -967 112560
rect -1289 108429 -967 108430
rect -1579 108302 -1452 108318
rect -1579 108178 -1475 108302
rect -1579 108162 -1452 108178
rect -2008 108050 -1686 108051
rect -2008 103920 -2007 108050
rect -1687 103920 -1686 108050
rect -2008 103919 -1686 103920
rect -2298 103792 -2171 103808
rect -2298 103668 -2194 103792
rect -2298 103652 -2171 103668
rect -2727 103540 -2405 103541
rect -2727 99410 -2726 103540
rect -2406 99410 -2405 103540
rect -2727 99409 -2405 99410
rect -2618 99031 -2514 99409
rect -2298 99298 -2251 103652
rect -2187 99298 -2171 103652
rect -1899 103541 -1795 103919
rect -1579 103808 -1532 108162
rect -1468 103808 -1452 108162
rect -1180 108051 -1076 108429
rect -860 108318 -813 112672
rect -749 108318 -733 112672
rect -461 112561 -357 112939
rect -141 112828 -94 117182
rect -30 112828 -14 117182
rect 258 117071 362 117449
rect 578 117338 625 121692
rect 689 117338 705 121692
rect 977 121581 1081 121959
rect 1297 121848 1344 126202
rect 1408 121848 1424 126202
rect 1696 126091 1800 126469
rect 2016 126358 2063 130712
rect 2127 126358 2143 130712
rect 2415 130601 2519 130979
rect 2735 130868 2782 135222
rect 2846 130868 2862 135222
rect 2735 130852 2862 130868
rect 2735 130728 2839 130852
rect 2735 130712 2862 130728
rect 2306 130600 2628 130601
rect 2306 126470 2307 130600
rect 2627 126470 2628 130600
rect 2306 126469 2628 126470
rect 2016 126342 2143 126358
rect 2016 126218 2120 126342
rect 2016 126202 2143 126218
rect 1587 126090 1909 126091
rect 1587 121960 1588 126090
rect 1908 121960 1909 126090
rect 1587 121959 1909 121960
rect 1297 121832 1424 121848
rect 1297 121708 1401 121832
rect 1297 121692 1424 121708
rect 868 121580 1190 121581
rect 868 117450 869 121580
rect 1189 117450 1190 121580
rect 868 117449 1190 117450
rect 578 117322 705 117338
rect 578 117198 682 117322
rect 578 117182 705 117198
rect 149 117070 471 117071
rect 149 112940 150 117070
rect 470 112940 471 117070
rect 149 112939 471 112940
rect -141 112812 -14 112828
rect -141 112688 -37 112812
rect -141 112672 -14 112688
rect -570 112560 -248 112561
rect -570 108430 -569 112560
rect -249 108430 -248 112560
rect -570 108429 -248 108430
rect -860 108302 -733 108318
rect -860 108178 -756 108302
rect -860 108162 -733 108178
rect -1289 108050 -967 108051
rect -1289 103920 -1288 108050
rect -968 103920 -967 108050
rect -1289 103919 -967 103920
rect -1579 103792 -1452 103808
rect -1579 103668 -1475 103792
rect -1579 103652 -1452 103668
rect -2008 103540 -1686 103541
rect -2008 99410 -2007 103540
rect -1687 99410 -1686 103540
rect -2008 99409 -1686 99410
rect -2298 99282 -2171 99298
rect -2298 99158 -2194 99282
rect -2298 99142 -2171 99158
rect -2727 99030 -2405 99031
rect -2727 94900 -2726 99030
rect -2406 94900 -2405 99030
rect -2727 94899 -2405 94900
rect -2618 94521 -2514 94899
rect -2298 94788 -2251 99142
rect -2187 94788 -2171 99142
rect -1899 99031 -1795 99409
rect -1579 99298 -1532 103652
rect -1468 99298 -1452 103652
rect -1180 103541 -1076 103919
rect -860 103808 -813 108162
rect -749 103808 -733 108162
rect -461 108051 -357 108429
rect -141 108318 -94 112672
rect -30 108318 -14 112672
rect 258 112561 362 112939
rect 578 112828 625 117182
rect 689 112828 705 117182
rect 977 117071 1081 117449
rect 1297 117338 1344 121692
rect 1408 117338 1424 121692
rect 1696 121581 1800 121959
rect 2016 121848 2063 126202
rect 2127 121848 2143 126202
rect 2415 126091 2519 126469
rect 2735 126358 2782 130712
rect 2846 126358 2862 130712
rect 2735 126342 2862 126358
rect 2735 126218 2839 126342
rect 2735 126202 2862 126218
rect 2306 126090 2628 126091
rect 2306 121960 2307 126090
rect 2627 121960 2628 126090
rect 2306 121959 2628 121960
rect 2016 121832 2143 121848
rect 2016 121708 2120 121832
rect 2016 121692 2143 121708
rect 1587 121580 1909 121581
rect 1587 117450 1588 121580
rect 1908 117450 1909 121580
rect 1587 117449 1909 117450
rect 1297 117322 1424 117338
rect 1297 117198 1401 117322
rect 1297 117182 1424 117198
rect 868 117070 1190 117071
rect 868 112940 869 117070
rect 1189 112940 1190 117070
rect 868 112939 1190 112940
rect 578 112812 705 112828
rect 578 112688 682 112812
rect 578 112672 705 112688
rect 149 112560 471 112561
rect 149 108430 150 112560
rect 470 108430 471 112560
rect 149 108429 471 108430
rect -141 108302 -14 108318
rect -141 108178 -37 108302
rect -141 108162 -14 108178
rect -570 108050 -248 108051
rect -570 103920 -569 108050
rect -249 103920 -248 108050
rect -570 103919 -248 103920
rect -860 103792 -733 103808
rect -860 103668 -756 103792
rect -860 103652 -733 103668
rect -1289 103540 -967 103541
rect -1289 99410 -1288 103540
rect -968 99410 -967 103540
rect -1289 99409 -967 99410
rect -1579 99282 -1452 99298
rect -1579 99158 -1475 99282
rect -1579 99142 -1452 99158
rect -2008 99030 -1686 99031
rect -2008 94900 -2007 99030
rect -1687 94900 -1686 99030
rect -2008 94899 -1686 94900
rect -2298 94772 -2171 94788
rect -2298 94648 -2194 94772
rect -2298 94632 -2171 94648
rect -2727 94520 -2405 94521
rect -2727 90390 -2726 94520
rect -2406 90390 -2405 94520
rect -2727 90389 -2405 90390
rect -2618 90011 -2514 90389
rect -2298 90278 -2251 94632
rect -2187 90278 -2171 94632
rect -1899 94521 -1795 94899
rect -1579 94788 -1532 99142
rect -1468 94788 -1452 99142
rect -1180 99031 -1076 99409
rect -860 99298 -813 103652
rect -749 99298 -733 103652
rect -461 103541 -357 103919
rect -141 103808 -94 108162
rect -30 103808 -14 108162
rect 258 108051 362 108429
rect 578 108318 625 112672
rect 689 108318 705 112672
rect 977 112561 1081 112939
rect 1297 112828 1344 117182
rect 1408 112828 1424 117182
rect 1696 117071 1800 117449
rect 2016 117338 2063 121692
rect 2127 117338 2143 121692
rect 2415 121581 2519 121959
rect 2735 121848 2782 126202
rect 2846 121848 2862 126202
rect 2735 121832 2862 121848
rect 2735 121708 2839 121832
rect 2735 121692 2862 121708
rect 2306 121580 2628 121581
rect 2306 117450 2307 121580
rect 2627 117450 2628 121580
rect 2306 117449 2628 117450
rect 2016 117322 2143 117338
rect 2016 117198 2120 117322
rect 2016 117182 2143 117198
rect 1587 117070 1909 117071
rect 1587 112940 1588 117070
rect 1908 112940 1909 117070
rect 1587 112939 1909 112940
rect 1297 112812 1424 112828
rect 1297 112688 1401 112812
rect 1297 112672 1424 112688
rect 868 112560 1190 112561
rect 868 108430 869 112560
rect 1189 108430 1190 112560
rect 868 108429 1190 108430
rect 578 108302 705 108318
rect 578 108178 682 108302
rect 578 108162 705 108178
rect 149 108050 471 108051
rect 149 103920 150 108050
rect 470 103920 471 108050
rect 149 103919 471 103920
rect -141 103792 -14 103808
rect -141 103668 -37 103792
rect -141 103652 -14 103668
rect -570 103540 -248 103541
rect -570 99410 -569 103540
rect -249 99410 -248 103540
rect -570 99409 -248 99410
rect -860 99282 -733 99298
rect -860 99158 -756 99282
rect -860 99142 -733 99158
rect -1289 99030 -967 99031
rect -1289 94900 -1288 99030
rect -968 94900 -967 99030
rect -1289 94899 -967 94900
rect -1579 94772 -1452 94788
rect -1579 94648 -1475 94772
rect -1579 94632 -1452 94648
rect -2008 94520 -1686 94521
rect -2008 90390 -2007 94520
rect -1687 90390 -1686 94520
rect -2008 90389 -1686 90390
rect -2298 90262 -2171 90278
rect -2298 90138 -2194 90262
rect -2298 90122 -2171 90138
rect -2727 90010 -2405 90011
rect -2727 85880 -2726 90010
rect -2406 85880 -2405 90010
rect -2727 85879 -2405 85880
rect -2618 85501 -2514 85879
rect -2298 85768 -2251 90122
rect -2187 85768 -2171 90122
rect -1899 90011 -1795 90389
rect -1579 90278 -1532 94632
rect -1468 90278 -1452 94632
rect -1180 94521 -1076 94899
rect -860 94788 -813 99142
rect -749 94788 -733 99142
rect -461 99031 -357 99409
rect -141 99298 -94 103652
rect -30 99298 -14 103652
rect 258 103541 362 103919
rect 578 103808 625 108162
rect 689 103808 705 108162
rect 977 108051 1081 108429
rect 1297 108318 1344 112672
rect 1408 108318 1424 112672
rect 1696 112561 1800 112939
rect 2016 112828 2063 117182
rect 2127 112828 2143 117182
rect 2415 117071 2519 117449
rect 2735 117338 2782 121692
rect 2846 117338 2862 121692
rect 2735 117322 2862 117338
rect 2735 117198 2839 117322
rect 2735 117182 2862 117198
rect 2306 117070 2628 117071
rect 2306 112940 2307 117070
rect 2627 112940 2628 117070
rect 2306 112939 2628 112940
rect 2016 112812 2143 112828
rect 2016 112688 2120 112812
rect 2016 112672 2143 112688
rect 1587 112560 1909 112561
rect 1587 108430 1588 112560
rect 1908 108430 1909 112560
rect 1587 108429 1909 108430
rect 1297 108302 1424 108318
rect 1297 108178 1401 108302
rect 1297 108162 1424 108178
rect 868 108050 1190 108051
rect 868 103920 869 108050
rect 1189 103920 1190 108050
rect 868 103919 1190 103920
rect 578 103792 705 103808
rect 578 103668 682 103792
rect 578 103652 705 103668
rect 149 103540 471 103541
rect 149 99410 150 103540
rect 470 99410 471 103540
rect 149 99409 471 99410
rect -141 99282 -14 99298
rect -141 99158 -37 99282
rect -141 99142 -14 99158
rect -570 99030 -248 99031
rect -570 94900 -569 99030
rect -249 94900 -248 99030
rect -570 94899 -248 94900
rect -860 94772 -733 94788
rect -860 94648 -756 94772
rect -860 94632 -733 94648
rect -1289 94520 -967 94521
rect -1289 90390 -1288 94520
rect -968 90390 -967 94520
rect -1289 90389 -967 90390
rect -1579 90262 -1452 90278
rect -1579 90138 -1475 90262
rect -1579 90122 -1452 90138
rect -2008 90010 -1686 90011
rect -2008 85880 -2007 90010
rect -1687 85880 -1686 90010
rect -2008 85879 -1686 85880
rect -2298 85752 -2171 85768
rect -2298 85628 -2194 85752
rect -2298 85612 -2171 85628
rect -2727 85500 -2405 85501
rect -2727 81370 -2726 85500
rect -2406 81370 -2405 85500
rect -2727 81369 -2405 81370
rect -2618 80991 -2514 81369
rect -2298 81258 -2251 85612
rect -2187 81258 -2171 85612
rect -1899 85501 -1795 85879
rect -1579 85768 -1532 90122
rect -1468 85768 -1452 90122
rect -1180 90011 -1076 90389
rect -860 90278 -813 94632
rect -749 90278 -733 94632
rect -461 94521 -357 94899
rect -141 94788 -94 99142
rect -30 94788 -14 99142
rect 258 99031 362 99409
rect 578 99298 625 103652
rect 689 99298 705 103652
rect 977 103541 1081 103919
rect 1297 103808 1344 108162
rect 1408 103808 1424 108162
rect 1696 108051 1800 108429
rect 2016 108318 2063 112672
rect 2127 108318 2143 112672
rect 2415 112561 2519 112939
rect 2735 112828 2782 117182
rect 2846 112828 2862 117182
rect 2735 112812 2862 112828
rect 2735 112688 2839 112812
rect 2735 112672 2862 112688
rect 2306 112560 2628 112561
rect 2306 108430 2307 112560
rect 2627 108430 2628 112560
rect 2306 108429 2628 108430
rect 2016 108302 2143 108318
rect 2016 108178 2120 108302
rect 2016 108162 2143 108178
rect 1587 108050 1909 108051
rect 1587 103920 1588 108050
rect 1908 103920 1909 108050
rect 1587 103919 1909 103920
rect 1297 103792 1424 103808
rect 1297 103668 1401 103792
rect 1297 103652 1424 103668
rect 868 103540 1190 103541
rect 868 99410 869 103540
rect 1189 99410 1190 103540
rect 868 99409 1190 99410
rect 578 99282 705 99298
rect 578 99158 682 99282
rect 578 99142 705 99158
rect 149 99030 471 99031
rect 149 94900 150 99030
rect 470 94900 471 99030
rect 149 94899 471 94900
rect -141 94772 -14 94788
rect -141 94648 -37 94772
rect -141 94632 -14 94648
rect -570 94520 -248 94521
rect -570 90390 -569 94520
rect -249 90390 -248 94520
rect -570 90389 -248 90390
rect -860 90262 -733 90278
rect -860 90138 -756 90262
rect -860 90122 -733 90138
rect -1289 90010 -967 90011
rect -1289 85880 -1288 90010
rect -968 85880 -967 90010
rect -1289 85879 -967 85880
rect -1579 85752 -1452 85768
rect -1579 85628 -1475 85752
rect -1579 85612 -1452 85628
rect -2008 85500 -1686 85501
rect -2008 81370 -2007 85500
rect -1687 81370 -1686 85500
rect -2008 81369 -1686 81370
rect -2298 81242 -2171 81258
rect -2298 81118 -2194 81242
rect -2298 81102 -2171 81118
rect -2727 80990 -2405 80991
rect -2727 76860 -2726 80990
rect -2406 76860 -2405 80990
rect -2727 76859 -2405 76860
rect -2618 76481 -2514 76859
rect -2298 76748 -2251 81102
rect -2187 76748 -2171 81102
rect -1899 80991 -1795 81369
rect -1579 81258 -1532 85612
rect -1468 81258 -1452 85612
rect -1180 85501 -1076 85879
rect -860 85768 -813 90122
rect -749 85768 -733 90122
rect -461 90011 -357 90389
rect -141 90278 -94 94632
rect -30 90278 -14 94632
rect 258 94521 362 94899
rect 578 94788 625 99142
rect 689 94788 705 99142
rect 977 99031 1081 99409
rect 1297 99298 1344 103652
rect 1408 99298 1424 103652
rect 1696 103541 1800 103919
rect 2016 103808 2063 108162
rect 2127 103808 2143 108162
rect 2415 108051 2519 108429
rect 2735 108318 2782 112672
rect 2846 108318 2862 112672
rect 2735 108302 2862 108318
rect 2735 108178 2839 108302
rect 2735 108162 2862 108178
rect 2306 108050 2628 108051
rect 2306 103920 2307 108050
rect 2627 103920 2628 108050
rect 2306 103919 2628 103920
rect 2016 103792 2143 103808
rect 2016 103668 2120 103792
rect 2016 103652 2143 103668
rect 1587 103540 1909 103541
rect 1587 99410 1588 103540
rect 1908 99410 1909 103540
rect 1587 99409 1909 99410
rect 1297 99282 1424 99298
rect 1297 99158 1401 99282
rect 1297 99142 1424 99158
rect 868 99030 1190 99031
rect 868 94900 869 99030
rect 1189 94900 1190 99030
rect 868 94899 1190 94900
rect 578 94772 705 94788
rect 578 94648 682 94772
rect 578 94632 705 94648
rect 149 94520 471 94521
rect 149 90390 150 94520
rect 470 90390 471 94520
rect 149 90389 471 90390
rect -141 90262 -14 90278
rect -141 90138 -37 90262
rect -141 90122 -14 90138
rect -570 90010 -248 90011
rect -570 85880 -569 90010
rect -249 85880 -248 90010
rect -570 85879 -248 85880
rect -860 85752 -733 85768
rect -860 85628 -756 85752
rect -860 85612 -733 85628
rect -1289 85500 -967 85501
rect -1289 81370 -1288 85500
rect -968 81370 -967 85500
rect -1289 81369 -967 81370
rect -1579 81242 -1452 81258
rect -1579 81118 -1475 81242
rect -1579 81102 -1452 81118
rect -2008 80990 -1686 80991
rect -2008 76860 -2007 80990
rect -1687 76860 -1686 80990
rect -2008 76859 -1686 76860
rect -2298 76732 -2171 76748
rect -2298 76608 -2194 76732
rect -2298 76592 -2171 76608
rect -2727 76480 -2405 76481
rect -2727 72350 -2726 76480
rect -2406 72350 -2405 76480
rect -2727 72349 -2405 72350
rect -2618 71971 -2514 72349
rect -2298 72238 -2251 76592
rect -2187 72238 -2171 76592
rect -1899 76481 -1795 76859
rect -1579 76748 -1532 81102
rect -1468 76748 -1452 81102
rect -1180 80991 -1076 81369
rect -860 81258 -813 85612
rect -749 81258 -733 85612
rect -461 85501 -357 85879
rect -141 85768 -94 90122
rect -30 85768 -14 90122
rect 258 90011 362 90389
rect 578 90278 625 94632
rect 689 90278 705 94632
rect 977 94521 1081 94899
rect 1297 94788 1344 99142
rect 1408 94788 1424 99142
rect 1696 99031 1800 99409
rect 2016 99298 2063 103652
rect 2127 99298 2143 103652
rect 2415 103541 2519 103919
rect 2735 103808 2782 108162
rect 2846 103808 2862 108162
rect 2735 103792 2862 103808
rect 2735 103668 2839 103792
rect 2735 103652 2862 103668
rect 2306 103540 2628 103541
rect 2306 99410 2307 103540
rect 2627 99410 2628 103540
rect 2306 99409 2628 99410
rect 2016 99282 2143 99298
rect 2016 99158 2120 99282
rect 2016 99142 2143 99158
rect 1587 99030 1909 99031
rect 1587 94900 1588 99030
rect 1908 94900 1909 99030
rect 1587 94899 1909 94900
rect 1297 94772 1424 94788
rect 1297 94648 1401 94772
rect 1297 94632 1424 94648
rect 868 94520 1190 94521
rect 868 90390 869 94520
rect 1189 90390 1190 94520
rect 868 90389 1190 90390
rect 578 90262 705 90278
rect 578 90138 682 90262
rect 578 90122 705 90138
rect 149 90010 471 90011
rect 149 85880 150 90010
rect 470 85880 471 90010
rect 149 85879 471 85880
rect -141 85752 -14 85768
rect -141 85628 -37 85752
rect -141 85612 -14 85628
rect -570 85500 -248 85501
rect -570 81370 -569 85500
rect -249 81370 -248 85500
rect -570 81369 -248 81370
rect -860 81242 -733 81258
rect -860 81118 -756 81242
rect -860 81102 -733 81118
rect -1289 80990 -967 80991
rect -1289 76860 -1288 80990
rect -968 76860 -967 80990
rect -1289 76859 -967 76860
rect -1579 76732 -1452 76748
rect -1579 76608 -1475 76732
rect -1579 76592 -1452 76608
rect -2008 76480 -1686 76481
rect -2008 72350 -2007 76480
rect -1687 72350 -1686 76480
rect -2008 72349 -1686 72350
rect -2298 72222 -2171 72238
rect -2298 72098 -2194 72222
rect -2298 72082 -2171 72098
rect -2727 71970 -2405 71971
rect -2727 67840 -2726 71970
rect -2406 67840 -2405 71970
rect -2727 67839 -2405 67840
rect -2618 67461 -2514 67839
rect -2298 67728 -2251 72082
rect -2187 67728 -2171 72082
rect -1899 71971 -1795 72349
rect -1579 72238 -1532 76592
rect -1468 72238 -1452 76592
rect -1180 76481 -1076 76859
rect -860 76748 -813 81102
rect -749 76748 -733 81102
rect -461 80991 -357 81369
rect -141 81258 -94 85612
rect -30 81258 -14 85612
rect 258 85501 362 85879
rect 578 85768 625 90122
rect 689 85768 705 90122
rect 977 90011 1081 90389
rect 1297 90278 1344 94632
rect 1408 90278 1424 94632
rect 1696 94521 1800 94899
rect 2016 94788 2063 99142
rect 2127 94788 2143 99142
rect 2415 99031 2519 99409
rect 2735 99298 2782 103652
rect 2846 99298 2862 103652
rect 2735 99282 2862 99298
rect 2735 99158 2839 99282
rect 2735 99142 2862 99158
rect 2306 99030 2628 99031
rect 2306 94900 2307 99030
rect 2627 94900 2628 99030
rect 2306 94899 2628 94900
rect 2016 94772 2143 94788
rect 2016 94648 2120 94772
rect 2016 94632 2143 94648
rect 1587 94520 1909 94521
rect 1587 90390 1588 94520
rect 1908 90390 1909 94520
rect 1587 90389 1909 90390
rect 1297 90262 1424 90278
rect 1297 90138 1401 90262
rect 1297 90122 1424 90138
rect 868 90010 1190 90011
rect 868 85880 869 90010
rect 1189 85880 1190 90010
rect 868 85879 1190 85880
rect 578 85752 705 85768
rect 578 85628 682 85752
rect 578 85612 705 85628
rect 149 85500 471 85501
rect 149 81370 150 85500
rect 470 81370 471 85500
rect 149 81369 471 81370
rect -141 81242 -14 81258
rect -141 81118 -37 81242
rect -141 81102 -14 81118
rect -570 80990 -248 80991
rect -570 76860 -569 80990
rect -249 76860 -248 80990
rect -570 76859 -248 76860
rect -860 76732 -733 76748
rect -860 76608 -756 76732
rect -860 76592 -733 76608
rect -1289 76480 -967 76481
rect -1289 72350 -1288 76480
rect -968 72350 -967 76480
rect -1289 72349 -967 72350
rect -1579 72222 -1452 72238
rect -1579 72098 -1475 72222
rect -1579 72082 -1452 72098
rect -2008 71970 -1686 71971
rect -2008 67840 -2007 71970
rect -1687 67840 -1686 71970
rect -2008 67839 -1686 67840
rect -2298 67712 -2171 67728
rect -2298 67588 -2194 67712
rect -2298 67572 -2171 67588
rect -2727 67460 -2405 67461
rect -2727 63330 -2726 67460
rect -2406 63330 -2405 67460
rect -2727 63329 -2405 63330
rect -2618 62951 -2514 63329
rect -2298 63218 -2251 67572
rect -2187 63218 -2171 67572
rect -1899 67461 -1795 67839
rect -1579 67728 -1532 72082
rect -1468 67728 -1452 72082
rect -1180 71971 -1076 72349
rect -860 72238 -813 76592
rect -749 72238 -733 76592
rect -461 76481 -357 76859
rect -141 76748 -94 81102
rect -30 76748 -14 81102
rect 258 80991 362 81369
rect 578 81258 625 85612
rect 689 81258 705 85612
rect 977 85501 1081 85879
rect 1297 85768 1344 90122
rect 1408 85768 1424 90122
rect 1696 90011 1800 90389
rect 2016 90278 2063 94632
rect 2127 90278 2143 94632
rect 2415 94521 2519 94899
rect 2735 94788 2782 99142
rect 2846 94788 2862 99142
rect 2735 94772 2862 94788
rect 2735 94648 2839 94772
rect 2735 94632 2862 94648
rect 2306 94520 2628 94521
rect 2306 90390 2307 94520
rect 2627 90390 2628 94520
rect 2306 90389 2628 90390
rect 2016 90262 2143 90278
rect 2016 90138 2120 90262
rect 2016 90122 2143 90138
rect 1587 90010 1909 90011
rect 1587 85880 1588 90010
rect 1908 85880 1909 90010
rect 1587 85879 1909 85880
rect 1297 85752 1424 85768
rect 1297 85628 1401 85752
rect 1297 85612 1424 85628
rect 868 85500 1190 85501
rect 868 81370 869 85500
rect 1189 81370 1190 85500
rect 868 81369 1190 81370
rect 578 81242 705 81258
rect 578 81118 682 81242
rect 578 81102 705 81118
rect 149 80990 471 80991
rect 149 76860 150 80990
rect 470 76860 471 80990
rect 149 76859 471 76860
rect -141 76732 -14 76748
rect -141 76608 -37 76732
rect -141 76592 -14 76608
rect -570 76480 -248 76481
rect -570 72350 -569 76480
rect -249 72350 -248 76480
rect -570 72349 -248 72350
rect -860 72222 -733 72238
rect -860 72098 -756 72222
rect -860 72082 -733 72098
rect -1289 71970 -967 71971
rect -1289 67840 -1288 71970
rect -968 67840 -967 71970
rect -1289 67839 -967 67840
rect -1579 67712 -1452 67728
rect -1579 67588 -1475 67712
rect -1579 67572 -1452 67588
rect -2008 67460 -1686 67461
rect -2008 63330 -2007 67460
rect -1687 63330 -1686 67460
rect -2008 63329 -1686 63330
rect -2298 63202 -2171 63218
rect -2298 63078 -2194 63202
rect -2298 63062 -2171 63078
rect -2727 62950 -2405 62951
rect -2727 58820 -2726 62950
rect -2406 58820 -2405 62950
rect -2727 58819 -2405 58820
rect -2618 58441 -2514 58819
rect -2298 58708 -2251 63062
rect -2187 58708 -2171 63062
rect -1899 62951 -1795 63329
rect -1579 63218 -1532 67572
rect -1468 63218 -1452 67572
rect -1180 67461 -1076 67839
rect -860 67728 -813 72082
rect -749 67728 -733 72082
rect -461 71971 -357 72349
rect -141 72238 -94 76592
rect -30 72238 -14 76592
rect 258 76481 362 76859
rect 578 76748 625 81102
rect 689 76748 705 81102
rect 977 80991 1081 81369
rect 1297 81258 1344 85612
rect 1408 81258 1424 85612
rect 1696 85501 1800 85879
rect 2016 85768 2063 90122
rect 2127 85768 2143 90122
rect 2415 90011 2519 90389
rect 2735 90278 2782 94632
rect 2846 90278 2862 94632
rect 2735 90262 2862 90278
rect 2735 90138 2839 90262
rect 2735 90122 2862 90138
rect 2306 90010 2628 90011
rect 2306 85880 2307 90010
rect 2627 85880 2628 90010
rect 2306 85879 2628 85880
rect 2016 85752 2143 85768
rect 2016 85628 2120 85752
rect 2016 85612 2143 85628
rect 1587 85500 1909 85501
rect 1587 81370 1588 85500
rect 1908 81370 1909 85500
rect 1587 81369 1909 81370
rect 1297 81242 1424 81258
rect 1297 81118 1401 81242
rect 1297 81102 1424 81118
rect 868 80990 1190 80991
rect 868 76860 869 80990
rect 1189 76860 1190 80990
rect 868 76859 1190 76860
rect 578 76732 705 76748
rect 578 76608 682 76732
rect 578 76592 705 76608
rect 149 76480 471 76481
rect 149 72350 150 76480
rect 470 72350 471 76480
rect 149 72349 471 72350
rect -141 72222 -14 72238
rect -141 72098 -37 72222
rect -141 72082 -14 72098
rect -570 71970 -248 71971
rect -570 67840 -569 71970
rect -249 67840 -248 71970
rect -570 67839 -248 67840
rect -860 67712 -733 67728
rect -860 67588 -756 67712
rect -860 67572 -733 67588
rect -1289 67460 -967 67461
rect -1289 63330 -1288 67460
rect -968 63330 -967 67460
rect -1289 63329 -967 63330
rect -1579 63202 -1452 63218
rect -1579 63078 -1475 63202
rect -1579 63062 -1452 63078
rect -2008 62950 -1686 62951
rect -2008 58820 -2007 62950
rect -1687 58820 -1686 62950
rect -2008 58819 -1686 58820
rect -2298 58692 -2171 58708
rect -2298 58568 -2194 58692
rect -2298 58552 -2171 58568
rect -2727 58440 -2405 58441
rect -2727 54310 -2726 58440
rect -2406 54310 -2405 58440
rect -2727 54309 -2405 54310
rect -2618 53931 -2514 54309
rect -2298 54198 -2251 58552
rect -2187 54198 -2171 58552
rect -1899 58441 -1795 58819
rect -1579 58708 -1532 63062
rect -1468 58708 -1452 63062
rect -1180 62951 -1076 63329
rect -860 63218 -813 67572
rect -749 63218 -733 67572
rect -461 67461 -357 67839
rect -141 67728 -94 72082
rect -30 67728 -14 72082
rect 258 71971 362 72349
rect 578 72238 625 76592
rect 689 72238 705 76592
rect 977 76481 1081 76859
rect 1297 76748 1344 81102
rect 1408 76748 1424 81102
rect 1696 80991 1800 81369
rect 2016 81258 2063 85612
rect 2127 81258 2143 85612
rect 2415 85501 2519 85879
rect 2735 85768 2782 90122
rect 2846 85768 2862 90122
rect 2735 85752 2862 85768
rect 2735 85628 2839 85752
rect 2735 85612 2862 85628
rect 2306 85500 2628 85501
rect 2306 81370 2307 85500
rect 2627 81370 2628 85500
rect 2306 81369 2628 81370
rect 2016 81242 2143 81258
rect 2016 81118 2120 81242
rect 2016 81102 2143 81118
rect 1587 80990 1909 80991
rect 1587 76860 1588 80990
rect 1908 76860 1909 80990
rect 1587 76859 1909 76860
rect 1297 76732 1424 76748
rect 1297 76608 1401 76732
rect 1297 76592 1424 76608
rect 868 76480 1190 76481
rect 868 72350 869 76480
rect 1189 72350 1190 76480
rect 868 72349 1190 72350
rect 578 72222 705 72238
rect 578 72098 682 72222
rect 578 72082 705 72098
rect 149 71970 471 71971
rect 149 67840 150 71970
rect 470 67840 471 71970
rect 149 67839 471 67840
rect -141 67712 -14 67728
rect -141 67588 -37 67712
rect -141 67572 -14 67588
rect -570 67460 -248 67461
rect -570 63330 -569 67460
rect -249 63330 -248 67460
rect -570 63329 -248 63330
rect -860 63202 -733 63218
rect -860 63078 -756 63202
rect -860 63062 -733 63078
rect -1289 62950 -967 62951
rect -1289 58820 -1288 62950
rect -968 58820 -967 62950
rect -1289 58819 -967 58820
rect -1579 58692 -1452 58708
rect -1579 58568 -1475 58692
rect -1579 58552 -1452 58568
rect -2008 58440 -1686 58441
rect -2008 54310 -2007 58440
rect -1687 54310 -1686 58440
rect -2008 54309 -1686 54310
rect -2298 54182 -2171 54198
rect -2298 54058 -2194 54182
rect -2298 54042 -2171 54058
rect -2727 53930 -2405 53931
rect -2727 49800 -2726 53930
rect -2406 49800 -2405 53930
rect -2727 49799 -2405 49800
rect -2618 49421 -2514 49799
rect -2298 49688 -2251 54042
rect -2187 49688 -2171 54042
rect -1899 53931 -1795 54309
rect -1579 54198 -1532 58552
rect -1468 54198 -1452 58552
rect -1180 58441 -1076 58819
rect -860 58708 -813 63062
rect -749 58708 -733 63062
rect -461 62951 -357 63329
rect -141 63218 -94 67572
rect -30 63218 -14 67572
rect 258 67461 362 67839
rect 578 67728 625 72082
rect 689 67728 705 72082
rect 977 71971 1081 72349
rect 1297 72238 1344 76592
rect 1408 72238 1424 76592
rect 1696 76481 1800 76859
rect 2016 76748 2063 81102
rect 2127 76748 2143 81102
rect 2415 80991 2519 81369
rect 2735 81258 2782 85612
rect 2846 81258 2862 85612
rect 2735 81242 2862 81258
rect 2735 81118 2839 81242
rect 2735 81102 2862 81118
rect 2306 80990 2628 80991
rect 2306 76860 2307 80990
rect 2627 76860 2628 80990
rect 2306 76859 2628 76860
rect 2016 76732 2143 76748
rect 2016 76608 2120 76732
rect 2016 76592 2143 76608
rect 1587 76480 1909 76481
rect 1587 72350 1588 76480
rect 1908 72350 1909 76480
rect 1587 72349 1909 72350
rect 1297 72222 1424 72238
rect 1297 72098 1401 72222
rect 1297 72082 1424 72098
rect 868 71970 1190 71971
rect 868 67840 869 71970
rect 1189 67840 1190 71970
rect 868 67839 1190 67840
rect 578 67712 705 67728
rect 578 67588 682 67712
rect 578 67572 705 67588
rect 149 67460 471 67461
rect 149 63330 150 67460
rect 470 63330 471 67460
rect 149 63329 471 63330
rect -141 63202 -14 63218
rect -141 63078 -37 63202
rect -141 63062 -14 63078
rect -570 62950 -248 62951
rect -570 58820 -569 62950
rect -249 58820 -248 62950
rect -570 58819 -248 58820
rect -860 58692 -733 58708
rect -860 58568 -756 58692
rect -860 58552 -733 58568
rect -1289 58440 -967 58441
rect -1289 54310 -1288 58440
rect -968 54310 -967 58440
rect -1289 54309 -967 54310
rect -1579 54182 -1452 54198
rect -1579 54058 -1475 54182
rect -1579 54042 -1452 54058
rect -2008 53930 -1686 53931
rect -2008 49800 -2007 53930
rect -1687 49800 -1686 53930
rect -2008 49799 -1686 49800
rect -2298 49672 -2171 49688
rect -2298 49548 -2194 49672
rect -2298 49532 -2171 49548
rect -2727 49420 -2405 49421
rect -2727 45290 -2726 49420
rect -2406 45290 -2405 49420
rect -2727 45289 -2405 45290
rect -2618 44911 -2514 45289
rect -2298 45178 -2251 49532
rect -2187 45178 -2171 49532
rect -1899 49421 -1795 49799
rect -1579 49688 -1532 54042
rect -1468 49688 -1452 54042
rect -1180 53931 -1076 54309
rect -860 54198 -813 58552
rect -749 54198 -733 58552
rect -461 58441 -357 58819
rect -141 58708 -94 63062
rect -30 58708 -14 63062
rect 258 62951 362 63329
rect 578 63218 625 67572
rect 689 63218 705 67572
rect 977 67461 1081 67839
rect 1297 67728 1344 72082
rect 1408 67728 1424 72082
rect 1696 71971 1800 72349
rect 2016 72238 2063 76592
rect 2127 72238 2143 76592
rect 2415 76481 2519 76859
rect 2735 76748 2782 81102
rect 2846 76748 2862 81102
rect 2735 76732 2862 76748
rect 2735 76608 2839 76732
rect 2735 76592 2862 76608
rect 2306 76480 2628 76481
rect 2306 72350 2307 76480
rect 2627 72350 2628 76480
rect 2306 72349 2628 72350
rect 2016 72222 2143 72238
rect 2016 72098 2120 72222
rect 2016 72082 2143 72098
rect 1587 71970 1909 71971
rect 1587 67840 1588 71970
rect 1908 67840 1909 71970
rect 1587 67839 1909 67840
rect 1297 67712 1424 67728
rect 1297 67588 1401 67712
rect 1297 67572 1424 67588
rect 868 67460 1190 67461
rect 868 63330 869 67460
rect 1189 63330 1190 67460
rect 868 63329 1190 63330
rect 578 63202 705 63218
rect 578 63078 682 63202
rect 578 63062 705 63078
rect 149 62950 471 62951
rect 149 58820 150 62950
rect 470 58820 471 62950
rect 149 58819 471 58820
rect -141 58692 -14 58708
rect -141 58568 -37 58692
rect -141 58552 -14 58568
rect -570 58440 -248 58441
rect -570 54310 -569 58440
rect -249 54310 -248 58440
rect -570 54309 -248 54310
rect -860 54182 -733 54198
rect -860 54058 -756 54182
rect -860 54042 -733 54058
rect -1289 53930 -967 53931
rect -1289 49800 -1288 53930
rect -968 49800 -967 53930
rect -1289 49799 -967 49800
rect -1579 49672 -1452 49688
rect -1579 49548 -1475 49672
rect -1579 49532 -1452 49548
rect -2008 49420 -1686 49421
rect -2008 45290 -2007 49420
rect -1687 45290 -1686 49420
rect -2008 45289 -1686 45290
rect -2298 45162 -2171 45178
rect -2298 45038 -2194 45162
rect -2298 45022 -2171 45038
rect -2727 44910 -2405 44911
rect -2727 40780 -2726 44910
rect -2406 40780 -2405 44910
rect -2727 40779 -2405 40780
rect -2618 40401 -2514 40779
rect -2298 40668 -2251 45022
rect -2187 40668 -2171 45022
rect -1899 44911 -1795 45289
rect -1579 45178 -1532 49532
rect -1468 45178 -1452 49532
rect -1180 49421 -1076 49799
rect -860 49688 -813 54042
rect -749 49688 -733 54042
rect -461 53931 -357 54309
rect -141 54198 -94 58552
rect -30 54198 -14 58552
rect 258 58441 362 58819
rect 578 58708 625 63062
rect 689 58708 705 63062
rect 977 62951 1081 63329
rect 1297 63218 1344 67572
rect 1408 63218 1424 67572
rect 1696 67461 1800 67839
rect 2016 67728 2063 72082
rect 2127 67728 2143 72082
rect 2415 71971 2519 72349
rect 2735 72238 2782 76592
rect 2846 72238 2862 76592
rect 2735 72222 2862 72238
rect 2735 72098 2839 72222
rect 2735 72082 2862 72098
rect 2306 71970 2628 71971
rect 2306 67840 2307 71970
rect 2627 67840 2628 71970
rect 2306 67839 2628 67840
rect 2016 67712 2143 67728
rect 2016 67588 2120 67712
rect 2016 67572 2143 67588
rect 1587 67460 1909 67461
rect 1587 63330 1588 67460
rect 1908 63330 1909 67460
rect 1587 63329 1909 63330
rect 1297 63202 1424 63218
rect 1297 63078 1401 63202
rect 1297 63062 1424 63078
rect 868 62950 1190 62951
rect 868 58820 869 62950
rect 1189 58820 1190 62950
rect 868 58819 1190 58820
rect 578 58692 705 58708
rect 578 58568 682 58692
rect 578 58552 705 58568
rect 149 58440 471 58441
rect 149 54310 150 58440
rect 470 54310 471 58440
rect 149 54309 471 54310
rect -141 54182 -14 54198
rect -141 54058 -37 54182
rect -141 54042 -14 54058
rect -570 53930 -248 53931
rect -570 49800 -569 53930
rect -249 49800 -248 53930
rect -570 49799 -248 49800
rect -860 49672 -733 49688
rect -860 49548 -756 49672
rect -860 49532 -733 49548
rect -1289 49420 -967 49421
rect -1289 45290 -1288 49420
rect -968 45290 -967 49420
rect -1289 45289 -967 45290
rect -1579 45162 -1452 45178
rect -1579 45038 -1475 45162
rect -1579 45022 -1452 45038
rect -2008 44910 -1686 44911
rect -2008 40780 -2007 44910
rect -1687 40780 -1686 44910
rect -2008 40779 -1686 40780
rect -2298 40652 -2171 40668
rect -2298 40528 -2194 40652
rect -2298 40512 -2171 40528
rect -2727 40400 -2405 40401
rect -2727 36270 -2726 40400
rect -2406 36270 -2405 40400
rect -2727 36269 -2405 36270
rect -2618 35891 -2514 36269
rect -2298 36158 -2251 40512
rect -2187 36158 -2171 40512
rect -1899 40401 -1795 40779
rect -1579 40668 -1532 45022
rect -1468 40668 -1452 45022
rect -1180 44911 -1076 45289
rect -860 45178 -813 49532
rect -749 45178 -733 49532
rect -461 49421 -357 49799
rect -141 49688 -94 54042
rect -30 49688 -14 54042
rect 258 53931 362 54309
rect 578 54198 625 58552
rect 689 54198 705 58552
rect 977 58441 1081 58819
rect 1297 58708 1344 63062
rect 1408 58708 1424 63062
rect 1696 62951 1800 63329
rect 2016 63218 2063 67572
rect 2127 63218 2143 67572
rect 2415 67461 2519 67839
rect 2735 67728 2782 72082
rect 2846 67728 2862 72082
rect 2735 67712 2862 67728
rect 2735 67588 2839 67712
rect 2735 67572 2862 67588
rect 2306 67460 2628 67461
rect 2306 63330 2307 67460
rect 2627 63330 2628 67460
rect 2306 63329 2628 63330
rect 2016 63202 2143 63218
rect 2016 63078 2120 63202
rect 2016 63062 2143 63078
rect 1587 62950 1909 62951
rect 1587 58820 1588 62950
rect 1908 58820 1909 62950
rect 1587 58819 1909 58820
rect 1297 58692 1424 58708
rect 1297 58568 1401 58692
rect 1297 58552 1424 58568
rect 868 58440 1190 58441
rect 868 54310 869 58440
rect 1189 54310 1190 58440
rect 868 54309 1190 54310
rect 578 54182 705 54198
rect 578 54058 682 54182
rect 578 54042 705 54058
rect 149 53930 471 53931
rect 149 49800 150 53930
rect 470 49800 471 53930
rect 149 49799 471 49800
rect -141 49672 -14 49688
rect -141 49548 -37 49672
rect -141 49532 -14 49548
rect -570 49420 -248 49421
rect -570 45290 -569 49420
rect -249 45290 -248 49420
rect -570 45289 -248 45290
rect -860 45162 -733 45178
rect -860 45038 -756 45162
rect -860 45022 -733 45038
rect -1289 44910 -967 44911
rect -1289 40780 -1288 44910
rect -968 40780 -967 44910
rect -1289 40779 -967 40780
rect -1579 40652 -1452 40668
rect -1579 40528 -1475 40652
rect -1579 40512 -1452 40528
rect -2008 40400 -1686 40401
rect -2008 36270 -2007 40400
rect -1687 36270 -1686 40400
rect -2008 36269 -1686 36270
rect -2298 36142 -2171 36158
rect -2298 36018 -2194 36142
rect -2298 36002 -2171 36018
rect -2727 35890 -2405 35891
rect -2727 31760 -2726 35890
rect -2406 31760 -2405 35890
rect -2727 31759 -2405 31760
rect -2618 31381 -2514 31759
rect -2298 31648 -2251 36002
rect -2187 31648 -2171 36002
rect -1899 35891 -1795 36269
rect -1579 36158 -1532 40512
rect -1468 36158 -1452 40512
rect -1180 40401 -1076 40779
rect -860 40668 -813 45022
rect -749 40668 -733 45022
rect -461 44911 -357 45289
rect -141 45178 -94 49532
rect -30 45178 -14 49532
rect 258 49421 362 49799
rect 578 49688 625 54042
rect 689 49688 705 54042
rect 977 53931 1081 54309
rect 1297 54198 1344 58552
rect 1408 54198 1424 58552
rect 1696 58441 1800 58819
rect 2016 58708 2063 63062
rect 2127 58708 2143 63062
rect 2415 62951 2519 63329
rect 2735 63218 2782 67572
rect 2846 63218 2862 67572
rect 2735 63202 2862 63218
rect 2735 63078 2839 63202
rect 2735 63062 2862 63078
rect 2306 62950 2628 62951
rect 2306 58820 2307 62950
rect 2627 58820 2628 62950
rect 2306 58819 2628 58820
rect 2016 58692 2143 58708
rect 2016 58568 2120 58692
rect 2016 58552 2143 58568
rect 1587 58440 1909 58441
rect 1587 54310 1588 58440
rect 1908 54310 1909 58440
rect 1587 54309 1909 54310
rect 1297 54182 1424 54198
rect 1297 54058 1401 54182
rect 1297 54042 1424 54058
rect 868 53930 1190 53931
rect 868 49800 869 53930
rect 1189 49800 1190 53930
rect 868 49799 1190 49800
rect 578 49672 705 49688
rect 578 49548 682 49672
rect 578 49532 705 49548
rect 149 49420 471 49421
rect 149 45290 150 49420
rect 470 45290 471 49420
rect 149 45289 471 45290
rect -141 45162 -14 45178
rect -141 45038 -37 45162
rect -141 45022 -14 45038
rect -570 44910 -248 44911
rect -570 40780 -569 44910
rect -249 40780 -248 44910
rect -570 40779 -248 40780
rect -860 40652 -733 40668
rect -860 40528 -756 40652
rect -860 40512 -733 40528
rect -1289 40400 -967 40401
rect -1289 36270 -1288 40400
rect -968 36270 -967 40400
rect -1289 36269 -967 36270
rect -1579 36142 -1452 36158
rect -1579 36018 -1475 36142
rect -1579 36002 -1452 36018
rect -2008 35890 -1686 35891
rect -2008 31760 -2007 35890
rect -1687 31760 -1686 35890
rect -2008 31759 -1686 31760
rect -2298 31632 -2171 31648
rect -2298 31508 -2194 31632
rect -2298 31492 -2171 31508
rect -2727 31380 -2405 31381
rect -2727 27250 -2726 31380
rect -2406 27250 -2405 31380
rect -2727 27249 -2405 27250
rect -2618 26871 -2514 27249
rect -2298 27138 -2251 31492
rect -2187 27138 -2171 31492
rect -1899 31381 -1795 31759
rect -1579 31648 -1532 36002
rect -1468 31648 -1452 36002
rect -1180 35891 -1076 36269
rect -860 36158 -813 40512
rect -749 36158 -733 40512
rect -461 40401 -357 40779
rect -141 40668 -94 45022
rect -30 40668 -14 45022
rect 258 44911 362 45289
rect 578 45178 625 49532
rect 689 45178 705 49532
rect 977 49421 1081 49799
rect 1297 49688 1344 54042
rect 1408 49688 1424 54042
rect 1696 53931 1800 54309
rect 2016 54198 2063 58552
rect 2127 54198 2143 58552
rect 2415 58441 2519 58819
rect 2735 58708 2782 63062
rect 2846 58708 2862 63062
rect 2735 58692 2862 58708
rect 2735 58568 2839 58692
rect 2735 58552 2862 58568
rect 2306 58440 2628 58441
rect 2306 54310 2307 58440
rect 2627 54310 2628 58440
rect 2306 54309 2628 54310
rect 2016 54182 2143 54198
rect 2016 54058 2120 54182
rect 2016 54042 2143 54058
rect 1587 53930 1909 53931
rect 1587 49800 1588 53930
rect 1908 49800 1909 53930
rect 1587 49799 1909 49800
rect 1297 49672 1424 49688
rect 1297 49548 1401 49672
rect 1297 49532 1424 49548
rect 868 49420 1190 49421
rect 868 45290 869 49420
rect 1189 45290 1190 49420
rect 868 45289 1190 45290
rect 578 45162 705 45178
rect 578 45038 682 45162
rect 578 45022 705 45038
rect 149 44910 471 44911
rect 149 40780 150 44910
rect 470 40780 471 44910
rect 149 40779 471 40780
rect -141 40652 -14 40668
rect -141 40528 -37 40652
rect -141 40512 -14 40528
rect -570 40400 -248 40401
rect -570 36270 -569 40400
rect -249 36270 -248 40400
rect -570 36269 -248 36270
rect -860 36142 -733 36158
rect -860 36018 -756 36142
rect -860 36002 -733 36018
rect -1289 35890 -967 35891
rect -1289 31760 -1288 35890
rect -968 31760 -967 35890
rect -1289 31759 -967 31760
rect -1579 31632 -1452 31648
rect -1579 31508 -1475 31632
rect -1579 31492 -1452 31508
rect -2008 31380 -1686 31381
rect -2008 27250 -2007 31380
rect -1687 27250 -1686 31380
rect -2008 27249 -1686 27250
rect -2298 27122 -2171 27138
rect -2298 26998 -2194 27122
rect -2298 26982 -2171 26998
rect -2727 26870 -2405 26871
rect -2727 22740 -2726 26870
rect -2406 22740 -2405 26870
rect -2727 22739 -2405 22740
rect -2618 22361 -2514 22739
rect -2298 22628 -2251 26982
rect -2187 22628 -2171 26982
rect -1899 26871 -1795 27249
rect -1579 27138 -1532 31492
rect -1468 27138 -1452 31492
rect -1180 31381 -1076 31759
rect -860 31648 -813 36002
rect -749 31648 -733 36002
rect -461 35891 -357 36269
rect -141 36158 -94 40512
rect -30 36158 -14 40512
rect 258 40401 362 40779
rect 578 40668 625 45022
rect 689 40668 705 45022
rect 977 44911 1081 45289
rect 1297 45178 1344 49532
rect 1408 45178 1424 49532
rect 1696 49421 1800 49799
rect 2016 49688 2063 54042
rect 2127 49688 2143 54042
rect 2415 53931 2519 54309
rect 2735 54198 2782 58552
rect 2846 54198 2862 58552
rect 2735 54182 2862 54198
rect 2735 54058 2839 54182
rect 2735 54042 2862 54058
rect 2306 53930 2628 53931
rect 2306 49800 2307 53930
rect 2627 49800 2628 53930
rect 2306 49799 2628 49800
rect 2016 49672 2143 49688
rect 2016 49548 2120 49672
rect 2016 49532 2143 49548
rect 1587 49420 1909 49421
rect 1587 45290 1588 49420
rect 1908 45290 1909 49420
rect 1587 45289 1909 45290
rect 1297 45162 1424 45178
rect 1297 45038 1401 45162
rect 1297 45022 1424 45038
rect 868 44910 1190 44911
rect 868 40780 869 44910
rect 1189 40780 1190 44910
rect 868 40779 1190 40780
rect 578 40652 705 40668
rect 578 40528 682 40652
rect 578 40512 705 40528
rect 149 40400 471 40401
rect 149 36270 150 40400
rect 470 36270 471 40400
rect 149 36269 471 36270
rect -141 36142 -14 36158
rect -141 36018 -37 36142
rect -141 36002 -14 36018
rect -570 35890 -248 35891
rect -570 31760 -569 35890
rect -249 31760 -248 35890
rect -570 31759 -248 31760
rect -860 31632 -733 31648
rect -860 31508 -756 31632
rect -860 31492 -733 31508
rect -1289 31380 -967 31381
rect -1289 27250 -1288 31380
rect -968 27250 -967 31380
rect -1289 27249 -967 27250
rect -1579 27122 -1452 27138
rect -1579 26998 -1475 27122
rect -1579 26982 -1452 26998
rect -2008 26870 -1686 26871
rect -2008 22740 -2007 26870
rect -1687 22740 -1686 26870
rect -2008 22739 -1686 22740
rect -2298 22612 -2171 22628
rect -2298 22488 -2194 22612
rect -2298 22472 -2171 22488
rect -2727 22360 -2405 22361
rect -2727 18230 -2726 22360
rect -2406 18230 -2405 22360
rect -2727 18229 -2405 18230
rect -2618 17851 -2514 18229
rect -2298 18118 -2251 22472
rect -2187 18118 -2171 22472
rect -1899 22361 -1795 22739
rect -1579 22628 -1532 26982
rect -1468 22628 -1452 26982
rect -1180 26871 -1076 27249
rect -860 27138 -813 31492
rect -749 27138 -733 31492
rect -461 31381 -357 31759
rect -141 31648 -94 36002
rect -30 31648 -14 36002
rect 258 35891 362 36269
rect 578 36158 625 40512
rect 689 36158 705 40512
rect 977 40401 1081 40779
rect 1297 40668 1344 45022
rect 1408 40668 1424 45022
rect 1696 44911 1800 45289
rect 2016 45178 2063 49532
rect 2127 45178 2143 49532
rect 2415 49421 2519 49799
rect 2735 49688 2782 54042
rect 2846 49688 2862 54042
rect 2735 49672 2862 49688
rect 2735 49548 2839 49672
rect 2735 49532 2862 49548
rect 2306 49420 2628 49421
rect 2306 45290 2307 49420
rect 2627 45290 2628 49420
rect 2306 45289 2628 45290
rect 2016 45162 2143 45178
rect 2016 45038 2120 45162
rect 2016 45022 2143 45038
rect 1587 44910 1909 44911
rect 1587 40780 1588 44910
rect 1908 40780 1909 44910
rect 1587 40779 1909 40780
rect 1297 40652 1424 40668
rect 1297 40528 1401 40652
rect 1297 40512 1424 40528
rect 868 40400 1190 40401
rect 868 36270 869 40400
rect 1189 36270 1190 40400
rect 868 36269 1190 36270
rect 578 36142 705 36158
rect 578 36018 682 36142
rect 578 36002 705 36018
rect 149 35890 471 35891
rect 149 31760 150 35890
rect 470 31760 471 35890
rect 149 31759 471 31760
rect -141 31632 -14 31648
rect -141 31508 -37 31632
rect -141 31492 -14 31508
rect -570 31380 -248 31381
rect -570 27250 -569 31380
rect -249 27250 -248 31380
rect -570 27249 -248 27250
rect -860 27122 -733 27138
rect -860 26998 -756 27122
rect -860 26982 -733 26998
rect -1289 26870 -967 26871
rect -1289 22740 -1288 26870
rect -968 22740 -967 26870
rect -1289 22739 -967 22740
rect -1579 22612 -1452 22628
rect -1579 22488 -1475 22612
rect -1579 22472 -1452 22488
rect -2008 22360 -1686 22361
rect -2008 18230 -2007 22360
rect -1687 18230 -1686 22360
rect -2008 18229 -1686 18230
rect -2298 18102 -2171 18118
rect -2298 17978 -2194 18102
rect -2298 17962 -2171 17978
rect -2727 17850 -2405 17851
rect -2727 13720 -2726 17850
rect -2406 13720 -2405 17850
rect -2727 13719 -2405 13720
rect -2618 13341 -2514 13719
rect -2298 13608 -2251 17962
rect -2187 13608 -2171 17962
rect -1899 17851 -1795 18229
rect -1579 18118 -1532 22472
rect -1468 18118 -1452 22472
rect -1180 22361 -1076 22739
rect -860 22628 -813 26982
rect -749 22628 -733 26982
rect -461 26871 -357 27249
rect -141 27138 -94 31492
rect -30 27138 -14 31492
rect 258 31381 362 31759
rect 578 31648 625 36002
rect 689 31648 705 36002
rect 977 35891 1081 36269
rect 1297 36158 1344 40512
rect 1408 36158 1424 40512
rect 1696 40401 1800 40779
rect 2016 40668 2063 45022
rect 2127 40668 2143 45022
rect 2415 44911 2519 45289
rect 2735 45178 2782 49532
rect 2846 45178 2862 49532
rect 2735 45162 2862 45178
rect 2735 45038 2839 45162
rect 2735 45022 2862 45038
rect 2306 44910 2628 44911
rect 2306 40780 2307 44910
rect 2627 40780 2628 44910
rect 2306 40779 2628 40780
rect 2016 40652 2143 40668
rect 2016 40528 2120 40652
rect 2016 40512 2143 40528
rect 1587 40400 1909 40401
rect 1587 36270 1588 40400
rect 1908 36270 1909 40400
rect 1587 36269 1909 36270
rect 1297 36142 1424 36158
rect 1297 36018 1401 36142
rect 1297 36002 1424 36018
rect 868 35890 1190 35891
rect 868 31760 869 35890
rect 1189 31760 1190 35890
rect 868 31759 1190 31760
rect 578 31632 705 31648
rect 578 31508 682 31632
rect 578 31492 705 31508
rect 149 31380 471 31381
rect 149 27250 150 31380
rect 470 27250 471 31380
rect 149 27249 471 27250
rect -141 27122 -14 27138
rect -141 26998 -37 27122
rect -141 26982 -14 26998
rect -570 26870 -248 26871
rect -570 22740 -569 26870
rect -249 22740 -248 26870
rect -570 22739 -248 22740
rect -860 22612 -733 22628
rect -860 22488 -756 22612
rect -860 22472 -733 22488
rect -1289 22360 -967 22361
rect -1289 18230 -1288 22360
rect -968 18230 -967 22360
rect -1289 18229 -967 18230
rect -1579 18102 -1452 18118
rect -1579 17978 -1475 18102
rect -1579 17962 -1452 17978
rect -2008 17850 -1686 17851
rect -2008 13720 -2007 17850
rect -1687 13720 -1686 17850
rect -2008 13719 -1686 13720
rect -2298 13592 -2171 13608
rect -2298 13468 -2194 13592
rect -2298 13452 -2171 13468
rect -2727 13340 -2405 13341
rect -2727 9210 -2726 13340
rect -2406 9210 -2405 13340
rect -2727 9209 -2405 9210
rect -2618 8831 -2514 9209
rect -2298 9098 -2251 13452
rect -2187 9098 -2171 13452
rect -1899 13341 -1795 13719
rect -1579 13608 -1532 17962
rect -1468 13608 -1452 17962
rect -1180 17851 -1076 18229
rect -860 18118 -813 22472
rect -749 18118 -733 22472
rect -461 22361 -357 22739
rect -141 22628 -94 26982
rect -30 22628 -14 26982
rect 258 26871 362 27249
rect 578 27138 625 31492
rect 689 27138 705 31492
rect 977 31381 1081 31759
rect 1297 31648 1344 36002
rect 1408 31648 1424 36002
rect 1696 35891 1800 36269
rect 2016 36158 2063 40512
rect 2127 36158 2143 40512
rect 2415 40401 2519 40779
rect 2735 40668 2782 45022
rect 2846 40668 2862 45022
rect 2735 40652 2862 40668
rect 2735 40528 2839 40652
rect 2735 40512 2862 40528
rect 2306 40400 2628 40401
rect 2306 36270 2307 40400
rect 2627 36270 2628 40400
rect 2306 36269 2628 36270
rect 2016 36142 2143 36158
rect 2016 36018 2120 36142
rect 2016 36002 2143 36018
rect 1587 35890 1909 35891
rect 1587 31760 1588 35890
rect 1908 31760 1909 35890
rect 1587 31759 1909 31760
rect 1297 31632 1424 31648
rect 1297 31508 1401 31632
rect 1297 31492 1424 31508
rect 868 31380 1190 31381
rect 868 27250 869 31380
rect 1189 27250 1190 31380
rect 868 27249 1190 27250
rect 578 27122 705 27138
rect 578 26998 682 27122
rect 578 26982 705 26998
rect 149 26870 471 26871
rect 149 22740 150 26870
rect 470 22740 471 26870
rect 149 22739 471 22740
rect -141 22612 -14 22628
rect -141 22488 -37 22612
rect -141 22472 -14 22488
rect -570 22360 -248 22361
rect -570 18230 -569 22360
rect -249 18230 -248 22360
rect -570 18229 -248 18230
rect -860 18102 -733 18118
rect -860 17978 -756 18102
rect -860 17962 -733 17978
rect -1289 17850 -967 17851
rect -1289 13720 -1288 17850
rect -968 13720 -967 17850
rect -1289 13719 -967 13720
rect -1579 13592 -1452 13608
rect -1579 13468 -1475 13592
rect -1579 13452 -1452 13468
rect -2008 13340 -1686 13341
rect -2008 9210 -2007 13340
rect -1687 9210 -1686 13340
rect -2008 9209 -1686 9210
rect -2298 9082 -2171 9098
rect -2298 8958 -2194 9082
rect -2298 8942 -2171 8958
rect -2727 8830 -2405 8831
rect -2727 4700 -2726 8830
rect -2406 4700 -2405 8830
rect -2727 4699 -2405 4700
rect -2618 4321 -2514 4699
rect -2298 4588 -2251 8942
rect -2187 4588 -2171 8942
rect -1899 8831 -1795 9209
rect -1579 9098 -1532 13452
rect -1468 9098 -1452 13452
rect -1180 13341 -1076 13719
rect -860 13608 -813 17962
rect -749 13608 -733 17962
rect -461 17851 -357 18229
rect -141 18118 -94 22472
rect -30 18118 -14 22472
rect 258 22361 362 22739
rect 578 22628 625 26982
rect 689 22628 705 26982
rect 977 26871 1081 27249
rect 1297 27138 1344 31492
rect 1408 27138 1424 31492
rect 1696 31381 1800 31759
rect 2016 31648 2063 36002
rect 2127 31648 2143 36002
rect 2415 35891 2519 36269
rect 2735 36158 2782 40512
rect 2846 36158 2862 40512
rect 2735 36142 2862 36158
rect 2735 36018 2839 36142
rect 2735 36002 2862 36018
rect 2306 35890 2628 35891
rect 2306 31760 2307 35890
rect 2627 31760 2628 35890
rect 2306 31759 2628 31760
rect 2016 31632 2143 31648
rect 2016 31508 2120 31632
rect 2016 31492 2143 31508
rect 1587 31380 1909 31381
rect 1587 27250 1588 31380
rect 1908 27250 1909 31380
rect 1587 27249 1909 27250
rect 1297 27122 1424 27138
rect 1297 26998 1401 27122
rect 1297 26982 1424 26998
rect 868 26870 1190 26871
rect 868 22740 869 26870
rect 1189 22740 1190 26870
rect 868 22739 1190 22740
rect 578 22612 705 22628
rect 578 22488 682 22612
rect 578 22472 705 22488
rect 149 22360 471 22361
rect 149 18230 150 22360
rect 470 18230 471 22360
rect 149 18229 471 18230
rect -141 18102 -14 18118
rect -141 17978 -37 18102
rect -141 17962 -14 17978
rect -570 17850 -248 17851
rect -570 13720 -569 17850
rect -249 13720 -248 17850
rect -570 13719 -248 13720
rect -860 13592 -733 13608
rect -860 13468 -756 13592
rect -860 13452 -733 13468
rect -1289 13340 -967 13341
rect -1289 9210 -1288 13340
rect -968 9210 -967 13340
rect -1289 9209 -967 9210
rect -1579 9082 -1452 9098
rect -1579 8958 -1475 9082
rect -1579 8942 -1452 8958
rect -2008 8830 -1686 8831
rect -2008 4700 -2007 8830
rect -1687 4700 -1686 8830
rect -2008 4699 -1686 4700
rect -2298 4572 -2171 4588
rect -2298 4448 -2194 4572
rect -2298 4432 -2171 4448
rect -2727 4320 -2405 4321
rect -2727 190 -2726 4320
rect -2406 190 -2405 4320
rect -2727 189 -2405 190
rect -2618 -189 -2514 189
rect -2298 78 -2251 4432
rect -2187 78 -2171 4432
rect -1899 4321 -1795 4699
rect -1579 4588 -1532 8942
rect -1468 4588 -1452 8942
rect -1180 8831 -1076 9209
rect -860 9098 -813 13452
rect -749 9098 -733 13452
rect -461 13341 -357 13719
rect -141 13608 -94 17962
rect -30 13608 -14 17962
rect 258 17851 362 18229
rect 578 18118 625 22472
rect 689 18118 705 22472
rect 977 22361 1081 22739
rect 1297 22628 1344 26982
rect 1408 22628 1424 26982
rect 1696 26871 1800 27249
rect 2016 27138 2063 31492
rect 2127 27138 2143 31492
rect 2415 31381 2519 31759
rect 2735 31648 2782 36002
rect 2846 31648 2862 36002
rect 2735 31632 2862 31648
rect 2735 31508 2839 31632
rect 2735 31492 2862 31508
rect 2306 31380 2628 31381
rect 2306 27250 2307 31380
rect 2627 27250 2628 31380
rect 2306 27249 2628 27250
rect 2016 27122 2143 27138
rect 2016 26998 2120 27122
rect 2016 26982 2143 26998
rect 1587 26870 1909 26871
rect 1587 22740 1588 26870
rect 1908 22740 1909 26870
rect 1587 22739 1909 22740
rect 1297 22612 1424 22628
rect 1297 22488 1401 22612
rect 1297 22472 1424 22488
rect 868 22360 1190 22361
rect 868 18230 869 22360
rect 1189 18230 1190 22360
rect 868 18229 1190 18230
rect 578 18102 705 18118
rect 578 17978 682 18102
rect 578 17962 705 17978
rect 149 17850 471 17851
rect 149 13720 150 17850
rect 470 13720 471 17850
rect 149 13719 471 13720
rect -141 13592 -14 13608
rect -141 13468 -37 13592
rect -141 13452 -14 13468
rect -570 13340 -248 13341
rect -570 9210 -569 13340
rect -249 9210 -248 13340
rect -570 9209 -248 9210
rect -860 9082 -733 9098
rect -860 8958 -756 9082
rect -860 8942 -733 8958
rect -1289 8830 -967 8831
rect -1289 4700 -1288 8830
rect -968 4700 -967 8830
rect -1289 4699 -967 4700
rect -1579 4572 -1452 4588
rect -1579 4448 -1475 4572
rect -1579 4432 -1452 4448
rect -2008 4320 -1686 4321
rect -2008 190 -2007 4320
rect -1687 190 -1686 4320
rect -2008 189 -1686 190
rect -2298 62 -2171 78
rect -2298 -62 -2194 62
rect -2298 -78 -2171 -62
rect -2727 -190 -2405 -189
rect -2727 -4320 -2726 -190
rect -2406 -4320 -2405 -190
rect -2727 -4321 -2405 -4320
rect -2618 -4699 -2514 -4321
rect -2298 -4432 -2251 -78
rect -2187 -4432 -2171 -78
rect -1899 -189 -1795 189
rect -1579 78 -1532 4432
rect -1468 78 -1452 4432
rect -1180 4321 -1076 4699
rect -860 4588 -813 8942
rect -749 4588 -733 8942
rect -461 8831 -357 9209
rect -141 9098 -94 13452
rect -30 9098 -14 13452
rect 258 13341 362 13719
rect 578 13608 625 17962
rect 689 13608 705 17962
rect 977 17851 1081 18229
rect 1297 18118 1344 22472
rect 1408 18118 1424 22472
rect 1696 22361 1800 22739
rect 2016 22628 2063 26982
rect 2127 22628 2143 26982
rect 2415 26871 2519 27249
rect 2735 27138 2782 31492
rect 2846 27138 2862 31492
rect 2735 27122 2862 27138
rect 2735 26998 2839 27122
rect 2735 26982 2862 26998
rect 2306 26870 2628 26871
rect 2306 22740 2307 26870
rect 2627 22740 2628 26870
rect 2306 22739 2628 22740
rect 2016 22612 2143 22628
rect 2016 22488 2120 22612
rect 2016 22472 2143 22488
rect 1587 22360 1909 22361
rect 1587 18230 1588 22360
rect 1908 18230 1909 22360
rect 1587 18229 1909 18230
rect 1297 18102 1424 18118
rect 1297 17978 1401 18102
rect 1297 17962 1424 17978
rect 868 17850 1190 17851
rect 868 13720 869 17850
rect 1189 13720 1190 17850
rect 868 13719 1190 13720
rect 578 13592 705 13608
rect 578 13468 682 13592
rect 578 13452 705 13468
rect 149 13340 471 13341
rect 149 9210 150 13340
rect 470 9210 471 13340
rect 149 9209 471 9210
rect -141 9082 -14 9098
rect -141 8958 -37 9082
rect -141 8942 -14 8958
rect -570 8830 -248 8831
rect -570 4700 -569 8830
rect -249 4700 -248 8830
rect -570 4699 -248 4700
rect -860 4572 -733 4588
rect -860 4448 -756 4572
rect -860 4432 -733 4448
rect -1289 4320 -967 4321
rect -1289 190 -1288 4320
rect -968 190 -967 4320
rect -1289 189 -967 190
rect -1579 62 -1452 78
rect -1579 -62 -1475 62
rect -1579 -78 -1452 -62
rect -2008 -190 -1686 -189
rect -2008 -4320 -2007 -190
rect -1687 -4320 -1686 -190
rect -2008 -4321 -1686 -4320
rect -2298 -4448 -2171 -4432
rect -2298 -4572 -2194 -4448
rect -2298 -4588 -2171 -4572
rect -2727 -4700 -2405 -4699
rect -2727 -8830 -2726 -4700
rect -2406 -8830 -2405 -4700
rect -2727 -8831 -2405 -8830
rect -2618 -9209 -2514 -8831
rect -2298 -8942 -2251 -4588
rect -2187 -8942 -2171 -4588
rect -1899 -4699 -1795 -4321
rect -1579 -4432 -1532 -78
rect -1468 -4432 -1452 -78
rect -1180 -189 -1076 189
rect -860 78 -813 4432
rect -749 78 -733 4432
rect -461 4321 -357 4699
rect -141 4588 -94 8942
rect -30 4588 -14 8942
rect 258 8831 362 9209
rect 578 9098 625 13452
rect 689 9098 705 13452
rect 977 13341 1081 13719
rect 1297 13608 1344 17962
rect 1408 13608 1424 17962
rect 1696 17851 1800 18229
rect 2016 18118 2063 22472
rect 2127 18118 2143 22472
rect 2415 22361 2519 22739
rect 2735 22628 2782 26982
rect 2846 22628 2862 26982
rect 2735 22612 2862 22628
rect 2735 22488 2839 22612
rect 2735 22472 2862 22488
rect 2306 22360 2628 22361
rect 2306 18230 2307 22360
rect 2627 18230 2628 22360
rect 2306 18229 2628 18230
rect 2016 18102 2143 18118
rect 2016 17978 2120 18102
rect 2016 17962 2143 17978
rect 1587 17850 1909 17851
rect 1587 13720 1588 17850
rect 1908 13720 1909 17850
rect 1587 13719 1909 13720
rect 1297 13592 1424 13608
rect 1297 13468 1401 13592
rect 1297 13452 1424 13468
rect 868 13340 1190 13341
rect 868 9210 869 13340
rect 1189 9210 1190 13340
rect 868 9209 1190 9210
rect 578 9082 705 9098
rect 578 8958 682 9082
rect 578 8942 705 8958
rect 149 8830 471 8831
rect 149 4700 150 8830
rect 470 4700 471 8830
rect 149 4699 471 4700
rect -141 4572 -14 4588
rect -141 4448 -37 4572
rect -141 4432 -14 4448
rect -570 4320 -248 4321
rect -570 190 -569 4320
rect -249 190 -248 4320
rect -570 189 -248 190
rect -860 62 -733 78
rect -860 -62 -756 62
rect -860 -78 -733 -62
rect -1289 -190 -967 -189
rect -1289 -4320 -1288 -190
rect -968 -4320 -967 -190
rect -1289 -4321 -967 -4320
rect -1579 -4448 -1452 -4432
rect -1579 -4572 -1475 -4448
rect -1579 -4588 -1452 -4572
rect -2008 -4700 -1686 -4699
rect -2008 -8830 -2007 -4700
rect -1687 -8830 -1686 -4700
rect -2008 -8831 -1686 -8830
rect -2298 -8958 -2171 -8942
rect -2298 -9082 -2194 -8958
rect -2298 -9098 -2171 -9082
rect -2727 -9210 -2405 -9209
rect -2727 -13340 -2726 -9210
rect -2406 -13340 -2405 -9210
rect -2727 -13341 -2405 -13340
rect -2618 -13719 -2514 -13341
rect -2298 -13452 -2251 -9098
rect -2187 -13452 -2171 -9098
rect -1899 -9209 -1795 -8831
rect -1579 -8942 -1532 -4588
rect -1468 -8942 -1452 -4588
rect -1180 -4699 -1076 -4321
rect -860 -4432 -813 -78
rect -749 -4432 -733 -78
rect -461 -189 -357 189
rect -141 78 -94 4432
rect -30 78 -14 4432
rect 258 4321 362 4699
rect 578 4588 625 8942
rect 689 4588 705 8942
rect 977 8831 1081 9209
rect 1297 9098 1344 13452
rect 1408 9098 1424 13452
rect 1696 13341 1800 13719
rect 2016 13608 2063 17962
rect 2127 13608 2143 17962
rect 2415 17851 2519 18229
rect 2735 18118 2782 22472
rect 2846 18118 2862 22472
rect 2735 18102 2862 18118
rect 2735 17978 2839 18102
rect 2735 17962 2862 17978
rect 2306 17850 2628 17851
rect 2306 13720 2307 17850
rect 2627 13720 2628 17850
rect 2306 13719 2628 13720
rect 2016 13592 2143 13608
rect 2016 13468 2120 13592
rect 2016 13452 2143 13468
rect 1587 13340 1909 13341
rect 1587 9210 1588 13340
rect 1908 9210 1909 13340
rect 1587 9209 1909 9210
rect 1297 9082 1424 9098
rect 1297 8958 1401 9082
rect 1297 8942 1424 8958
rect 868 8830 1190 8831
rect 868 4700 869 8830
rect 1189 4700 1190 8830
rect 868 4699 1190 4700
rect 578 4572 705 4588
rect 578 4448 682 4572
rect 578 4432 705 4448
rect 149 4320 471 4321
rect 149 190 150 4320
rect 470 190 471 4320
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -4320 -569 -190
rect -249 -4320 -248 -190
rect -570 -4321 -248 -4320
rect -860 -4448 -733 -4432
rect -860 -4572 -756 -4448
rect -860 -4588 -733 -4572
rect -1289 -4700 -967 -4699
rect -1289 -8830 -1288 -4700
rect -968 -8830 -967 -4700
rect -1289 -8831 -967 -8830
rect -1579 -8958 -1452 -8942
rect -1579 -9082 -1475 -8958
rect -1579 -9098 -1452 -9082
rect -2008 -9210 -1686 -9209
rect -2008 -13340 -2007 -9210
rect -1687 -13340 -1686 -9210
rect -2008 -13341 -1686 -13340
rect -2298 -13468 -2171 -13452
rect -2298 -13592 -2194 -13468
rect -2298 -13608 -2171 -13592
rect -2727 -13720 -2405 -13719
rect -2727 -17850 -2726 -13720
rect -2406 -17850 -2405 -13720
rect -2727 -17851 -2405 -17850
rect -2618 -18229 -2514 -17851
rect -2298 -17962 -2251 -13608
rect -2187 -17962 -2171 -13608
rect -1899 -13719 -1795 -13341
rect -1579 -13452 -1532 -9098
rect -1468 -13452 -1452 -9098
rect -1180 -9209 -1076 -8831
rect -860 -8942 -813 -4588
rect -749 -8942 -733 -4588
rect -461 -4699 -357 -4321
rect -141 -4432 -94 -78
rect -30 -4432 -14 -78
rect 258 -189 362 189
rect 578 78 625 4432
rect 689 78 705 4432
rect 977 4321 1081 4699
rect 1297 4588 1344 8942
rect 1408 4588 1424 8942
rect 1696 8831 1800 9209
rect 2016 9098 2063 13452
rect 2127 9098 2143 13452
rect 2415 13341 2519 13719
rect 2735 13608 2782 17962
rect 2846 13608 2862 17962
rect 2735 13592 2862 13608
rect 2735 13468 2839 13592
rect 2735 13452 2862 13468
rect 2306 13340 2628 13341
rect 2306 9210 2307 13340
rect 2627 9210 2628 13340
rect 2306 9209 2628 9210
rect 2016 9082 2143 9098
rect 2016 8958 2120 9082
rect 2016 8942 2143 8958
rect 1587 8830 1909 8831
rect 1587 4700 1588 8830
rect 1908 4700 1909 8830
rect 1587 4699 1909 4700
rect 1297 4572 1424 4588
rect 1297 4448 1401 4572
rect 1297 4432 1424 4448
rect 868 4320 1190 4321
rect 868 190 869 4320
rect 1189 190 1190 4320
rect 868 189 1190 190
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -4320 150 -190
rect 470 -4320 471 -190
rect 149 -4321 471 -4320
rect -141 -4448 -14 -4432
rect -141 -4572 -37 -4448
rect -141 -4588 -14 -4572
rect -570 -4700 -248 -4699
rect -570 -8830 -569 -4700
rect -249 -8830 -248 -4700
rect -570 -8831 -248 -8830
rect -860 -8958 -733 -8942
rect -860 -9082 -756 -8958
rect -860 -9098 -733 -9082
rect -1289 -9210 -967 -9209
rect -1289 -13340 -1288 -9210
rect -968 -13340 -967 -9210
rect -1289 -13341 -967 -13340
rect -1579 -13468 -1452 -13452
rect -1579 -13592 -1475 -13468
rect -1579 -13608 -1452 -13592
rect -2008 -13720 -1686 -13719
rect -2008 -17850 -2007 -13720
rect -1687 -17850 -1686 -13720
rect -2008 -17851 -1686 -17850
rect -2298 -17978 -2171 -17962
rect -2298 -18102 -2194 -17978
rect -2298 -18118 -2171 -18102
rect -2727 -18230 -2405 -18229
rect -2727 -22360 -2726 -18230
rect -2406 -22360 -2405 -18230
rect -2727 -22361 -2405 -22360
rect -2618 -22739 -2514 -22361
rect -2298 -22472 -2251 -18118
rect -2187 -22472 -2171 -18118
rect -1899 -18229 -1795 -17851
rect -1579 -17962 -1532 -13608
rect -1468 -17962 -1452 -13608
rect -1180 -13719 -1076 -13341
rect -860 -13452 -813 -9098
rect -749 -13452 -733 -9098
rect -461 -9209 -357 -8831
rect -141 -8942 -94 -4588
rect -30 -8942 -14 -4588
rect 258 -4699 362 -4321
rect 578 -4432 625 -78
rect 689 -4432 705 -78
rect 977 -189 1081 189
rect 1297 78 1344 4432
rect 1408 78 1424 4432
rect 1696 4321 1800 4699
rect 2016 4588 2063 8942
rect 2127 4588 2143 8942
rect 2415 8831 2519 9209
rect 2735 9098 2782 13452
rect 2846 9098 2862 13452
rect 2735 9082 2862 9098
rect 2735 8958 2839 9082
rect 2735 8942 2862 8958
rect 2306 8830 2628 8831
rect 2306 4700 2307 8830
rect 2627 4700 2628 8830
rect 2306 4699 2628 4700
rect 2016 4572 2143 4588
rect 2016 4448 2120 4572
rect 2016 4432 2143 4448
rect 1587 4320 1909 4321
rect 1587 190 1588 4320
rect 1908 190 1909 4320
rect 1587 189 1909 190
rect 1297 62 1424 78
rect 1297 -62 1401 62
rect 1297 -78 1424 -62
rect 868 -190 1190 -189
rect 868 -4320 869 -190
rect 1189 -4320 1190 -190
rect 868 -4321 1190 -4320
rect 578 -4448 705 -4432
rect 578 -4572 682 -4448
rect 578 -4588 705 -4572
rect 149 -4700 471 -4699
rect 149 -8830 150 -4700
rect 470 -8830 471 -4700
rect 149 -8831 471 -8830
rect -141 -8958 -14 -8942
rect -141 -9082 -37 -8958
rect -141 -9098 -14 -9082
rect -570 -9210 -248 -9209
rect -570 -13340 -569 -9210
rect -249 -13340 -248 -9210
rect -570 -13341 -248 -13340
rect -860 -13468 -733 -13452
rect -860 -13592 -756 -13468
rect -860 -13608 -733 -13592
rect -1289 -13720 -967 -13719
rect -1289 -17850 -1288 -13720
rect -968 -17850 -967 -13720
rect -1289 -17851 -967 -17850
rect -1579 -17978 -1452 -17962
rect -1579 -18102 -1475 -17978
rect -1579 -18118 -1452 -18102
rect -2008 -18230 -1686 -18229
rect -2008 -22360 -2007 -18230
rect -1687 -22360 -1686 -18230
rect -2008 -22361 -1686 -22360
rect -2298 -22488 -2171 -22472
rect -2298 -22612 -2194 -22488
rect -2298 -22628 -2171 -22612
rect -2727 -22740 -2405 -22739
rect -2727 -26870 -2726 -22740
rect -2406 -26870 -2405 -22740
rect -2727 -26871 -2405 -26870
rect -2618 -27249 -2514 -26871
rect -2298 -26982 -2251 -22628
rect -2187 -26982 -2171 -22628
rect -1899 -22739 -1795 -22361
rect -1579 -22472 -1532 -18118
rect -1468 -22472 -1452 -18118
rect -1180 -18229 -1076 -17851
rect -860 -17962 -813 -13608
rect -749 -17962 -733 -13608
rect -461 -13719 -357 -13341
rect -141 -13452 -94 -9098
rect -30 -13452 -14 -9098
rect 258 -9209 362 -8831
rect 578 -8942 625 -4588
rect 689 -8942 705 -4588
rect 977 -4699 1081 -4321
rect 1297 -4432 1344 -78
rect 1408 -4432 1424 -78
rect 1696 -189 1800 189
rect 2016 78 2063 4432
rect 2127 78 2143 4432
rect 2415 4321 2519 4699
rect 2735 4588 2782 8942
rect 2846 4588 2862 8942
rect 2735 4572 2862 4588
rect 2735 4448 2839 4572
rect 2735 4432 2862 4448
rect 2306 4320 2628 4321
rect 2306 190 2307 4320
rect 2627 190 2628 4320
rect 2306 189 2628 190
rect 2016 62 2143 78
rect 2016 -62 2120 62
rect 2016 -78 2143 -62
rect 1587 -190 1909 -189
rect 1587 -4320 1588 -190
rect 1908 -4320 1909 -190
rect 1587 -4321 1909 -4320
rect 1297 -4448 1424 -4432
rect 1297 -4572 1401 -4448
rect 1297 -4588 1424 -4572
rect 868 -4700 1190 -4699
rect 868 -8830 869 -4700
rect 1189 -8830 1190 -4700
rect 868 -8831 1190 -8830
rect 578 -8958 705 -8942
rect 578 -9082 682 -8958
rect 578 -9098 705 -9082
rect 149 -9210 471 -9209
rect 149 -13340 150 -9210
rect 470 -13340 471 -9210
rect 149 -13341 471 -13340
rect -141 -13468 -14 -13452
rect -141 -13592 -37 -13468
rect -141 -13608 -14 -13592
rect -570 -13720 -248 -13719
rect -570 -17850 -569 -13720
rect -249 -17850 -248 -13720
rect -570 -17851 -248 -17850
rect -860 -17978 -733 -17962
rect -860 -18102 -756 -17978
rect -860 -18118 -733 -18102
rect -1289 -18230 -967 -18229
rect -1289 -22360 -1288 -18230
rect -968 -22360 -967 -18230
rect -1289 -22361 -967 -22360
rect -1579 -22488 -1452 -22472
rect -1579 -22612 -1475 -22488
rect -1579 -22628 -1452 -22612
rect -2008 -22740 -1686 -22739
rect -2008 -26870 -2007 -22740
rect -1687 -26870 -1686 -22740
rect -2008 -26871 -1686 -26870
rect -2298 -26998 -2171 -26982
rect -2298 -27122 -2194 -26998
rect -2298 -27138 -2171 -27122
rect -2727 -27250 -2405 -27249
rect -2727 -31380 -2726 -27250
rect -2406 -31380 -2405 -27250
rect -2727 -31381 -2405 -31380
rect -2618 -31759 -2514 -31381
rect -2298 -31492 -2251 -27138
rect -2187 -31492 -2171 -27138
rect -1899 -27249 -1795 -26871
rect -1579 -26982 -1532 -22628
rect -1468 -26982 -1452 -22628
rect -1180 -22739 -1076 -22361
rect -860 -22472 -813 -18118
rect -749 -22472 -733 -18118
rect -461 -18229 -357 -17851
rect -141 -17962 -94 -13608
rect -30 -17962 -14 -13608
rect 258 -13719 362 -13341
rect 578 -13452 625 -9098
rect 689 -13452 705 -9098
rect 977 -9209 1081 -8831
rect 1297 -8942 1344 -4588
rect 1408 -8942 1424 -4588
rect 1696 -4699 1800 -4321
rect 2016 -4432 2063 -78
rect 2127 -4432 2143 -78
rect 2415 -189 2519 189
rect 2735 78 2782 4432
rect 2846 78 2862 4432
rect 2735 62 2862 78
rect 2735 -62 2839 62
rect 2735 -78 2862 -62
rect 2306 -190 2628 -189
rect 2306 -4320 2307 -190
rect 2627 -4320 2628 -190
rect 2306 -4321 2628 -4320
rect 2016 -4448 2143 -4432
rect 2016 -4572 2120 -4448
rect 2016 -4588 2143 -4572
rect 1587 -4700 1909 -4699
rect 1587 -8830 1588 -4700
rect 1908 -8830 1909 -4700
rect 1587 -8831 1909 -8830
rect 1297 -8958 1424 -8942
rect 1297 -9082 1401 -8958
rect 1297 -9098 1424 -9082
rect 868 -9210 1190 -9209
rect 868 -13340 869 -9210
rect 1189 -13340 1190 -9210
rect 868 -13341 1190 -13340
rect 578 -13468 705 -13452
rect 578 -13592 682 -13468
rect 578 -13608 705 -13592
rect 149 -13720 471 -13719
rect 149 -17850 150 -13720
rect 470 -17850 471 -13720
rect 149 -17851 471 -17850
rect -141 -17978 -14 -17962
rect -141 -18102 -37 -17978
rect -141 -18118 -14 -18102
rect -570 -18230 -248 -18229
rect -570 -22360 -569 -18230
rect -249 -22360 -248 -18230
rect -570 -22361 -248 -22360
rect -860 -22488 -733 -22472
rect -860 -22612 -756 -22488
rect -860 -22628 -733 -22612
rect -1289 -22740 -967 -22739
rect -1289 -26870 -1288 -22740
rect -968 -26870 -967 -22740
rect -1289 -26871 -967 -26870
rect -1579 -26998 -1452 -26982
rect -1579 -27122 -1475 -26998
rect -1579 -27138 -1452 -27122
rect -2008 -27250 -1686 -27249
rect -2008 -31380 -2007 -27250
rect -1687 -31380 -1686 -27250
rect -2008 -31381 -1686 -31380
rect -2298 -31508 -2171 -31492
rect -2298 -31632 -2194 -31508
rect -2298 -31648 -2171 -31632
rect -2727 -31760 -2405 -31759
rect -2727 -35890 -2726 -31760
rect -2406 -35890 -2405 -31760
rect -2727 -35891 -2405 -35890
rect -2618 -36269 -2514 -35891
rect -2298 -36002 -2251 -31648
rect -2187 -36002 -2171 -31648
rect -1899 -31759 -1795 -31381
rect -1579 -31492 -1532 -27138
rect -1468 -31492 -1452 -27138
rect -1180 -27249 -1076 -26871
rect -860 -26982 -813 -22628
rect -749 -26982 -733 -22628
rect -461 -22739 -357 -22361
rect -141 -22472 -94 -18118
rect -30 -22472 -14 -18118
rect 258 -18229 362 -17851
rect 578 -17962 625 -13608
rect 689 -17962 705 -13608
rect 977 -13719 1081 -13341
rect 1297 -13452 1344 -9098
rect 1408 -13452 1424 -9098
rect 1696 -9209 1800 -8831
rect 2016 -8942 2063 -4588
rect 2127 -8942 2143 -4588
rect 2415 -4699 2519 -4321
rect 2735 -4432 2782 -78
rect 2846 -4432 2862 -78
rect 2735 -4448 2862 -4432
rect 2735 -4572 2839 -4448
rect 2735 -4588 2862 -4572
rect 2306 -4700 2628 -4699
rect 2306 -8830 2307 -4700
rect 2627 -8830 2628 -4700
rect 2306 -8831 2628 -8830
rect 2016 -8958 2143 -8942
rect 2016 -9082 2120 -8958
rect 2016 -9098 2143 -9082
rect 1587 -9210 1909 -9209
rect 1587 -13340 1588 -9210
rect 1908 -13340 1909 -9210
rect 1587 -13341 1909 -13340
rect 1297 -13468 1424 -13452
rect 1297 -13592 1401 -13468
rect 1297 -13608 1424 -13592
rect 868 -13720 1190 -13719
rect 868 -17850 869 -13720
rect 1189 -17850 1190 -13720
rect 868 -17851 1190 -17850
rect 578 -17978 705 -17962
rect 578 -18102 682 -17978
rect 578 -18118 705 -18102
rect 149 -18230 471 -18229
rect 149 -22360 150 -18230
rect 470 -22360 471 -18230
rect 149 -22361 471 -22360
rect -141 -22488 -14 -22472
rect -141 -22612 -37 -22488
rect -141 -22628 -14 -22612
rect -570 -22740 -248 -22739
rect -570 -26870 -569 -22740
rect -249 -26870 -248 -22740
rect -570 -26871 -248 -26870
rect -860 -26998 -733 -26982
rect -860 -27122 -756 -26998
rect -860 -27138 -733 -27122
rect -1289 -27250 -967 -27249
rect -1289 -31380 -1288 -27250
rect -968 -31380 -967 -27250
rect -1289 -31381 -967 -31380
rect -1579 -31508 -1452 -31492
rect -1579 -31632 -1475 -31508
rect -1579 -31648 -1452 -31632
rect -2008 -31760 -1686 -31759
rect -2008 -35890 -2007 -31760
rect -1687 -35890 -1686 -31760
rect -2008 -35891 -1686 -35890
rect -2298 -36018 -2171 -36002
rect -2298 -36142 -2194 -36018
rect -2298 -36158 -2171 -36142
rect -2727 -36270 -2405 -36269
rect -2727 -40400 -2726 -36270
rect -2406 -40400 -2405 -36270
rect -2727 -40401 -2405 -40400
rect -2618 -40779 -2514 -40401
rect -2298 -40512 -2251 -36158
rect -2187 -40512 -2171 -36158
rect -1899 -36269 -1795 -35891
rect -1579 -36002 -1532 -31648
rect -1468 -36002 -1452 -31648
rect -1180 -31759 -1076 -31381
rect -860 -31492 -813 -27138
rect -749 -31492 -733 -27138
rect -461 -27249 -357 -26871
rect -141 -26982 -94 -22628
rect -30 -26982 -14 -22628
rect 258 -22739 362 -22361
rect 578 -22472 625 -18118
rect 689 -22472 705 -18118
rect 977 -18229 1081 -17851
rect 1297 -17962 1344 -13608
rect 1408 -17962 1424 -13608
rect 1696 -13719 1800 -13341
rect 2016 -13452 2063 -9098
rect 2127 -13452 2143 -9098
rect 2415 -9209 2519 -8831
rect 2735 -8942 2782 -4588
rect 2846 -8942 2862 -4588
rect 2735 -8958 2862 -8942
rect 2735 -9082 2839 -8958
rect 2735 -9098 2862 -9082
rect 2306 -9210 2628 -9209
rect 2306 -13340 2307 -9210
rect 2627 -13340 2628 -9210
rect 2306 -13341 2628 -13340
rect 2016 -13468 2143 -13452
rect 2016 -13592 2120 -13468
rect 2016 -13608 2143 -13592
rect 1587 -13720 1909 -13719
rect 1587 -17850 1588 -13720
rect 1908 -17850 1909 -13720
rect 1587 -17851 1909 -17850
rect 1297 -17978 1424 -17962
rect 1297 -18102 1401 -17978
rect 1297 -18118 1424 -18102
rect 868 -18230 1190 -18229
rect 868 -22360 869 -18230
rect 1189 -22360 1190 -18230
rect 868 -22361 1190 -22360
rect 578 -22488 705 -22472
rect 578 -22612 682 -22488
rect 578 -22628 705 -22612
rect 149 -22740 471 -22739
rect 149 -26870 150 -22740
rect 470 -26870 471 -22740
rect 149 -26871 471 -26870
rect -141 -26998 -14 -26982
rect -141 -27122 -37 -26998
rect -141 -27138 -14 -27122
rect -570 -27250 -248 -27249
rect -570 -31380 -569 -27250
rect -249 -31380 -248 -27250
rect -570 -31381 -248 -31380
rect -860 -31508 -733 -31492
rect -860 -31632 -756 -31508
rect -860 -31648 -733 -31632
rect -1289 -31760 -967 -31759
rect -1289 -35890 -1288 -31760
rect -968 -35890 -967 -31760
rect -1289 -35891 -967 -35890
rect -1579 -36018 -1452 -36002
rect -1579 -36142 -1475 -36018
rect -1579 -36158 -1452 -36142
rect -2008 -36270 -1686 -36269
rect -2008 -40400 -2007 -36270
rect -1687 -40400 -1686 -36270
rect -2008 -40401 -1686 -40400
rect -2298 -40528 -2171 -40512
rect -2298 -40652 -2194 -40528
rect -2298 -40668 -2171 -40652
rect -2727 -40780 -2405 -40779
rect -2727 -44910 -2726 -40780
rect -2406 -44910 -2405 -40780
rect -2727 -44911 -2405 -44910
rect -2618 -45289 -2514 -44911
rect -2298 -45022 -2251 -40668
rect -2187 -45022 -2171 -40668
rect -1899 -40779 -1795 -40401
rect -1579 -40512 -1532 -36158
rect -1468 -40512 -1452 -36158
rect -1180 -36269 -1076 -35891
rect -860 -36002 -813 -31648
rect -749 -36002 -733 -31648
rect -461 -31759 -357 -31381
rect -141 -31492 -94 -27138
rect -30 -31492 -14 -27138
rect 258 -27249 362 -26871
rect 578 -26982 625 -22628
rect 689 -26982 705 -22628
rect 977 -22739 1081 -22361
rect 1297 -22472 1344 -18118
rect 1408 -22472 1424 -18118
rect 1696 -18229 1800 -17851
rect 2016 -17962 2063 -13608
rect 2127 -17962 2143 -13608
rect 2415 -13719 2519 -13341
rect 2735 -13452 2782 -9098
rect 2846 -13452 2862 -9098
rect 2735 -13468 2862 -13452
rect 2735 -13592 2839 -13468
rect 2735 -13608 2862 -13592
rect 2306 -13720 2628 -13719
rect 2306 -17850 2307 -13720
rect 2627 -17850 2628 -13720
rect 2306 -17851 2628 -17850
rect 2016 -17978 2143 -17962
rect 2016 -18102 2120 -17978
rect 2016 -18118 2143 -18102
rect 1587 -18230 1909 -18229
rect 1587 -22360 1588 -18230
rect 1908 -22360 1909 -18230
rect 1587 -22361 1909 -22360
rect 1297 -22488 1424 -22472
rect 1297 -22612 1401 -22488
rect 1297 -22628 1424 -22612
rect 868 -22740 1190 -22739
rect 868 -26870 869 -22740
rect 1189 -26870 1190 -22740
rect 868 -26871 1190 -26870
rect 578 -26998 705 -26982
rect 578 -27122 682 -26998
rect 578 -27138 705 -27122
rect 149 -27250 471 -27249
rect 149 -31380 150 -27250
rect 470 -31380 471 -27250
rect 149 -31381 471 -31380
rect -141 -31508 -14 -31492
rect -141 -31632 -37 -31508
rect -141 -31648 -14 -31632
rect -570 -31760 -248 -31759
rect -570 -35890 -569 -31760
rect -249 -35890 -248 -31760
rect -570 -35891 -248 -35890
rect -860 -36018 -733 -36002
rect -860 -36142 -756 -36018
rect -860 -36158 -733 -36142
rect -1289 -36270 -967 -36269
rect -1289 -40400 -1288 -36270
rect -968 -40400 -967 -36270
rect -1289 -40401 -967 -40400
rect -1579 -40528 -1452 -40512
rect -1579 -40652 -1475 -40528
rect -1579 -40668 -1452 -40652
rect -2008 -40780 -1686 -40779
rect -2008 -44910 -2007 -40780
rect -1687 -44910 -1686 -40780
rect -2008 -44911 -1686 -44910
rect -2298 -45038 -2171 -45022
rect -2298 -45162 -2194 -45038
rect -2298 -45178 -2171 -45162
rect -2727 -45290 -2405 -45289
rect -2727 -49420 -2726 -45290
rect -2406 -49420 -2405 -45290
rect -2727 -49421 -2405 -49420
rect -2618 -49799 -2514 -49421
rect -2298 -49532 -2251 -45178
rect -2187 -49532 -2171 -45178
rect -1899 -45289 -1795 -44911
rect -1579 -45022 -1532 -40668
rect -1468 -45022 -1452 -40668
rect -1180 -40779 -1076 -40401
rect -860 -40512 -813 -36158
rect -749 -40512 -733 -36158
rect -461 -36269 -357 -35891
rect -141 -36002 -94 -31648
rect -30 -36002 -14 -31648
rect 258 -31759 362 -31381
rect 578 -31492 625 -27138
rect 689 -31492 705 -27138
rect 977 -27249 1081 -26871
rect 1297 -26982 1344 -22628
rect 1408 -26982 1424 -22628
rect 1696 -22739 1800 -22361
rect 2016 -22472 2063 -18118
rect 2127 -22472 2143 -18118
rect 2415 -18229 2519 -17851
rect 2735 -17962 2782 -13608
rect 2846 -17962 2862 -13608
rect 2735 -17978 2862 -17962
rect 2735 -18102 2839 -17978
rect 2735 -18118 2862 -18102
rect 2306 -18230 2628 -18229
rect 2306 -22360 2307 -18230
rect 2627 -22360 2628 -18230
rect 2306 -22361 2628 -22360
rect 2016 -22488 2143 -22472
rect 2016 -22612 2120 -22488
rect 2016 -22628 2143 -22612
rect 1587 -22740 1909 -22739
rect 1587 -26870 1588 -22740
rect 1908 -26870 1909 -22740
rect 1587 -26871 1909 -26870
rect 1297 -26998 1424 -26982
rect 1297 -27122 1401 -26998
rect 1297 -27138 1424 -27122
rect 868 -27250 1190 -27249
rect 868 -31380 869 -27250
rect 1189 -31380 1190 -27250
rect 868 -31381 1190 -31380
rect 578 -31508 705 -31492
rect 578 -31632 682 -31508
rect 578 -31648 705 -31632
rect 149 -31760 471 -31759
rect 149 -35890 150 -31760
rect 470 -35890 471 -31760
rect 149 -35891 471 -35890
rect -141 -36018 -14 -36002
rect -141 -36142 -37 -36018
rect -141 -36158 -14 -36142
rect -570 -36270 -248 -36269
rect -570 -40400 -569 -36270
rect -249 -40400 -248 -36270
rect -570 -40401 -248 -40400
rect -860 -40528 -733 -40512
rect -860 -40652 -756 -40528
rect -860 -40668 -733 -40652
rect -1289 -40780 -967 -40779
rect -1289 -44910 -1288 -40780
rect -968 -44910 -967 -40780
rect -1289 -44911 -967 -44910
rect -1579 -45038 -1452 -45022
rect -1579 -45162 -1475 -45038
rect -1579 -45178 -1452 -45162
rect -2008 -45290 -1686 -45289
rect -2008 -49420 -2007 -45290
rect -1687 -49420 -1686 -45290
rect -2008 -49421 -1686 -49420
rect -2298 -49548 -2171 -49532
rect -2298 -49672 -2194 -49548
rect -2298 -49688 -2171 -49672
rect -2727 -49800 -2405 -49799
rect -2727 -53930 -2726 -49800
rect -2406 -53930 -2405 -49800
rect -2727 -53931 -2405 -53930
rect -2618 -54309 -2514 -53931
rect -2298 -54042 -2251 -49688
rect -2187 -54042 -2171 -49688
rect -1899 -49799 -1795 -49421
rect -1579 -49532 -1532 -45178
rect -1468 -49532 -1452 -45178
rect -1180 -45289 -1076 -44911
rect -860 -45022 -813 -40668
rect -749 -45022 -733 -40668
rect -461 -40779 -357 -40401
rect -141 -40512 -94 -36158
rect -30 -40512 -14 -36158
rect 258 -36269 362 -35891
rect 578 -36002 625 -31648
rect 689 -36002 705 -31648
rect 977 -31759 1081 -31381
rect 1297 -31492 1344 -27138
rect 1408 -31492 1424 -27138
rect 1696 -27249 1800 -26871
rect 2016 -26982 2063 -22628
rect 2127 -26982 2143 -22628
rect 2415 -22739 2519 -22361
rect 2735 -22472 2782 -18118
rect 2846 -22472 2862 -18118
rect 2735 -22488 2862 -22472
rect 2735 -22612 2839 -22488
rect 2735 -22628 2862 -22612
rect 2306 -22740 2628 -22739
rect 2306 -26870 2307 -22740
rect 2627 -26870 2628 -22740
rect 2306 -26871 2628 -26870
rect 2016 -26998 2143 -26982
rect 2016 -27122 2120 -26998
rect 2016 -27138 2143 -27122
rect 1587 -27250 1909 -27249
rect 1587 -31380 1588 -27250
rect 1908 -31380 1909 -27250
rect 1587 -31381 1909 -31380
rect 1297 -31508 1424 -31492
rect 1297 -31632 1401 -31508
rect 1297 -31648 1424 -31632
rect 868 -31760 1190 -31759
rect 868 -35890 869 -31760
rect 1189 -35890 1190 -31760
rect 868 -35891 1190 -35890
rect 578 -36018 705 -36002
rect 578 -36142 682 -36018
rect 578 -36158 705 -36142
rect 149 -36270 471 -36269
rect 149 -40400 150 -36270
rect 470 -40400 471 -36270
rect 149 -40401 471 -40400
rect -141 -40528 -14 -40512
rect -141 -40652 -37 -40528
rect -141 -40668 -14 -40652
rect -570 -40780 -248 -40779
rect -570 -44910 -569 -40780
rect -249 -44910 -248 -40780
rect -570 -44911 -248 -44910
rect -860 -45038 -733 -45022
rect -860 -45162 -756 -45038
rect -860 -45178 -733 -45162
rect -1289 -45290 -967 -45289
rect -1289 -49420 -1288 -45290
rect -968 -49420 -967 -45290
rect -1289 -49421 -967 -49420
rect -1579 -49548 -1452 -49532
rect -1579 -49672 -1475 -49548
rect -1579 -49688 -1452 -49672
rect -2008 -49800 -1686 -49799
rect -2008 -53930 -2007 -49800
rect -1687 -53930 -1686 -49800
rect -2008 -53931 -1686 -53930
rect -2298 -54058 -2171 -54042
rect -2298 -54182 -2194 -54058
rect -2298 -54198 -2171 -54182
rect -2727 -54310 -2405 -54309
rect -2727 -58440 -2726 -54310
rect -2406 -58440 -2405 -54310
rect -2727 -58441 -2405 -58440
rect -2618 -58819 -2514 -58441
rect -2298 -58552 -2251 -54198
rect -2187 -58552 -2171 -54198
rect -1899 -54309 -1795 -53931
rect -1579 -54042 -1532 -49688
rect -1468 -54042 -1452 -49688
rect -1180 -49799 -1076 -49421
rect -860 -49532 -813 -45178
rect -749 -49532 -733 -45178
rect -461 -45289 -357 -44911
rect -141 -45022 -94 -40668
rect -30 -45022 -14 -40668
rect 258 -40779 362 -40401
rect 578 -40512 625 -36158
rect 689 -40512 705 -36158
rect 977 -36269 1081 -35891
rect 1297 -36002 1344 -31648
rect 1408 -36002 1424 -31648
rect 1696 -31759 1800 -31381
rect 2016 -31492 2063 -27138
rect 2127 -31492 2143 -27138
rect 2415 -27249 2519 -26871
rect 2735 -26982 2782 -22628
rect 2846 -26982 2862 -22628
rect 2735 -26998 2862 -26982
rect 2735 -27122 2839 -26998
rect 2735 -27138 2862 -27122
rect 2306 -27250 2628 -27249
rect 2306 -31380 2307 -27250
rect 2627 -31380 2628 -27250
rect 2306 -31381 2628 -31380
rect 2016 -31508 2143 -31492
rect 2016 -31632 2120 -31508
rect 2016 -31648 2143 -31632
rect 1587 -31760 1909 -31759
rect 1587 -35890 1588 -31760
rect 1908 -35890 1909 -31760
rect 1587 -35891 1909 -35890
rect 1297 -36018 1424 -36002
rect 1297 -36142 1401 -36018
rect 1297 -36158 1424 -36142
rect 868 -36270 1190 -36269
rect 868 -40400 869 -36270
rect 1189 -40400 1190 -36270
rect 868 -40401 1190 -40400
rect 578 -40528 705 -40512
rect 578 -40652 682 -40528
rect 578 -40668 705 -40652
rect 149 -40780 471 -40779
rect 149 -44910 150 -40780
rect 470 -44910 471 -40780
rect 149 -44911 471 -44910
rect -141 -45038 -14 -45022
rect -141 -45162 -37 -45038
rect -141 -45178 -14 -45162
rect -570 -45290 -248 -45289
rect -570 -49420 -569 -45290
rect -249 -49420 -248 -45290
rect -570 -49421 -248 -49420
rect -860 -49548 -733 -49532
rect -860 -49672 -756 -49548
rect -860 -49688 -733 -49672
rect -1289 -49800 -967 -49799
rect -1289 -53930 -1288 -49800
rect -968 -53930 -967 -49800
rect -1289 -53931 -967 -53930
rect -1579 -54058 -1452 -54042
rect -1579 -54182 -1475 -54058
rect -1579 -54198 -1452 -54182
rect -2008 -54310 -1686 -54309
rect -2008 -58440 -2007 -54310
rect -1687 -58440 -1686 -54310
rect -2008 -58441 -1686 -58440
rect -2298 -58568 -2171 -58552
rect -2298 -58692 -2194 -58568
rect -2298 -58708 -2171 -58692
rect -2727 -58820 -2405 -58819
rect -2727 -62950 -2726 -58820
rect -2406 -62950 -2405 -58820
rect -2727 -62951 -2405 -62950
rect -2618 -63329 -2514 -62951
rect -2298 -63062 -2251 -58708
rect -2187 -63062 -2171 -58708
rect -1899 -58819 -1795 -58441
rect -1579 -58552 -1532 -54198
rect -1468 -58552 -1452 -54198
rect -1180 -54309 -1076 -53931
rect -860 -54042 -813 -49688
rect -749 -54042 -733 -49688
rect -461 -49799 -357 -49421
rect -141 -49532 -94 -45178
rect -30 -49532 -14 -45178
rect 258 -45289 362 -44911
rect 578 -45022 625 -40668
rect 689 -45022 705 -40668
rect 977 -40779 1081 -40401
rect 1297 -40512 1344 -36158
rect 1408 -40512 1424 -36158
rect 1696 -36269 1800 -35891
rect 2016 -36002 2063 -31648
rect 2127 -36002 2143 -31648
rect 2415 -31759 2519 -31381
rect 2735 -31492 2782 -27138
rect 2846 -31492 2862 -27138
rect 2735 -31508 2862 -31492
rect 2735 -31632 2839 -31508
rect 2735 -31648 2862 -31632
rect 2306 -31760 2628 -31759
rect 2306 -35890 2307 -31760
rect 2627 -35890 2628 -31760
rect 2306 -35891 2628 -35890
rect 2016 -36018 2143 -36002
rect 2016 -36142 2120 -36018
rect 2016 -36158 2143 -36142
rect 1587 -36270 1909 -36269
rect 1587 -40400 1588 -36270
rect 1908 -40400 1909 -36270
rect 1587 -40401 1909 -40400
rect 1297 -40528 1424 -40512
rect 1297 -40652 1401 -40528
rect 1297 -40668 1424 -40652
rect 868 -40780 1190 -40779
rect 868 -44910 869 -40780
rect 1189 -44910 1190 -40780
rect 868 -44911 1190 -44910
rect 578 -45038 705 -45022
rect 578 -45162 682 -45038
rect 578 -45178 705 -45162
rect 149 -45290 471 -45289
rect 149 -49420 150 -45290
rect 470 -49420 471 -45290
rect 149 -49421 471 -49420
rect -141 -49548 -14 -49532
rect -141 -49672 -37 -49548
rect -141 -49688 -14 -49672
rect -570 -49800 -248 -49799
rect -570 -53930 -569 -49800
rect -249 -53930 -248 -49800
rect -570 -53931 -248 -53930
rect -860 -54058 -733 -54042
rect -860 -54182 -756 -54058
rect -860 -54198 -733 -54182
rect -1289 -54310 -967 -54309
rect -1289 -58440 -1288 -54310
rect -968 -58440 -967 -54310
rect -1289 -58441 -967 -58440
rect -1579 -58568 -1452 -58552
rect -1579 -58692 -1475 -58568
rect -1579 -58708 -1452 -58692
rect -2008 -58820 -1686 -58819
rect -2008 -62950 -2007 -58820
rect -1687 -62950 -1686 -58820
rect -2008 -62951 -1686 -62950
rect -2298 -63078 -2171 -63062
rect -2298 -63202 -2194 -63078
rect -2298 -63218 -2171 -63202
rect -2727 -63330 -2405 -63329
rect -2727 -67460 -2726 -63330
rect -2406 -67460 -2405 -63330
rect -2727 -67461 -2405 -67460
rect -2618 -67839 -2514 -67461
rect -2298 -67572 -2251 -63218
rect -2187 -67572 -2171 -63218
rect -1899 -63329 -1795 -62951
rect -1579 -63062 -1532 -58708
rect -1468 -63062 -1452 -58708
rect -1180 -58819 -1076 -58441
rect -860 -58552 -813 -54198
rect -749 -58552 -733 -54198
rect -461 -54309 -357 -53931
rect -141 -54042 -94 -49688
rect -30 -54042 -14 -49688
rect 258 -49799 362 -49421
rect 578 -49532 625 -45178
rect 689 -49532 705 -45178
rect 977 -45289 1081 -44911
rect 1297 -45022 1344 -40668
rect 1408 -45022 1424 -40668
rect 1696 -40779 1800 -40401
rect 2016 -40512 2063 -36158
rect 2127 -40512 2143 -36158
rect 2415 -36269 2519 -35891
rect 2735 -36002 2782 -31648
rect 2846 -36002 2862 -31648
rect 2735 -36018 2862 -36002
rect 2735 -36142 2839 -36018
rect 2735 -36158 2862 -36142
rect 2306 -36270 2628 -36269
rect 2306 -40400 2307 -36270
rect 2627 -40400 2628 -36270
rect 2306 -40401 2628 -40400
rect 2016 -40528 2143 -40512
rect 2016 -40652 2120 -40528
rect 2016 -40668 2143 -40652
rect 1587 -40780 1909 -40779
rect 1587 -44910 1588 -40780
rect 1908 -44910 1909 -40780
rect 1587 -44911 1909 -44910
rect 1297 -45038 1424 -45022
rect 1297 -45162 1401 -45038
rect 1297 -45178 1424 -45162
rect 868 -45290 1190 -45289
rect 868 -49420 869 -45290
rect 1189 -49420 1190 -45290
rect 868 -49421 1190 -49420
rect 578 -49548 705 -49532
rect 578 -49672 682 -49548
rect 578 -49688 705 -49672
rect 149 -49800 471 -49799
rect 149 -53930 150 -49800
rect 470 -53930 471 -49800
rect 149 -53931 471 -53930
rect -141 -54058 -14 -54042
rect -141 -54182 -37 -54058
rect -141 -54198 -14 -54182
rect -570 -54310 -248 -54309
rect -570 -58440 -569 -54310
rect -249 -58440 -248 -54310
rect -570 -58441 -248 -58440
rect -860 -58568 -733 -58552
rect -860 -58692 -756 -58568
rect -860 -58708 -733 -58692
rect -1289 -58820 -967 -58819
rect -1289 -62950 -1288 -58820
rect -968 -62950 -967 -58820
rect -1289 -62951 -967 -62950
rect -1579 -63078 -1452 -63062
rect -1579 -63202 -1475 -63078
rect -1579 -63218 -1452 -63202
rect -2008 -63330 -1686 -63329
rect -2008 -67460 -2007 -63330
rect -1687 -67460 -1686 -63330
rect -2008 -67461 -1686 -67460
rect -2298 -67588 -2171 -67572
rect -2298 -67712 -2194 -67588
rect -2298 -67728 -2171 -67712
rect -2727 -67840 -2405 -67839
rect -2727 -71970 -2726 -67840
rect -2406 -71970 -2405 -67840
rect -2727 -71971 -2405 -71970
rect -2618 -72349 -2514 -71971
rect -2298 -72082 -2251 -67728
rect -2187 -72082 -2171 -67728
rect -1899 -67839 -1795 -67461
rect -1579 -67572 -1532 -63218
rect -1468 -67572 -1452 -63218
rect -1180 -63329 -1076 -62951
rect -860 -63062 -813 -58708
rect -749 -63062 -733 -58708
rect -461 -58819 -357 -58441
rect -141 -58552 -94 -54198
rect -30 -58552 -14 -54198
rect 258 -54309 362 -53931
rect 578 -54042 625 -49688
rect 689 -54042 705 -49688
rect 977 -49799 1081 -49421
rect 1297 -49532 1344 -45178
rect 1408 -49532 1424 -45178
rect 1696 -45289 1800 -44911
rect 2016 -45022 2063 -40668
rect 2127 -45022 2143 -40668
rect 2415 -40779 2519 -40401
rect 2735 -40512 2782 -36158
rect 2846 -40512 2862 -36158
rect 2735 -40528 2862 -40512
rect 2735 -40652 2839 -40528
rect 2735 -40668 2862 -40652
rect 2306 -40780 2628 -40779
rect 2306 -44910 2307 -40780
rect 2627 -44910 2628 -40780
rect 2306 -44911 2628 -44910
rect 2016 -45038 2143 -45022
rect 2016 -45162 2120 -45038
rect 2016 -45178 2143 -45162
rect 1587 -45290 1909 -45289
rect 1587 -49420 1588 -45290
rect 1908 -49420 1909 -45290
rect 1587 -49421 1909 -49420
rect 1297 -49548 1424 -49532
rect 1297 -49672 1401 -49548
rect 1297 -49688 1424 -49672
rect 868 -49800 1190 -49799
rect 868 -53930 869 -49800
rect 1189 -53930 1190 -49800
rect 868 -53931 1190 -53930
rect 578 -54058 705 -54042
rect 578 -54182 682 -54058
rect 578 -54198 705 -54182
rect 149 -54310 471 -54309
rect 149 -58440 150 -54310
rect 470 -58440 471 -54310
rect 149 -58441 471 -58440
rect -141 -58568 -14 -58552
rect -141 -58692 -37 -58568
rect -141 -58708 -14 -58692
rect -570 -58820 -248 -58819
rect -570 -62950 -569 -58820
rect -249 -62950 -248 -58820
rect -570 -62951 -248 -62950
rect -860 -63078 -733 -63062
rect -860 -63202 -756 -63078
rect -860 -63218 -733 -63202
rect -1289 -63330 -967 -63329
rect -1289 -67460 -1288 -63330
rect -968 -67460 -967 -63330
rect -1289 -67461 -967 -67460
rect -1579 -67588 -1452 -67572
rect -1579 -67712 -1475 -67588
rect -1579 -67728 -1452 -67712
rect -2008 -67840 -1686 -67839
rect -2008 -71970 -2007 -67840
rect -1687 -71970 -1686 -67840
rect -2008 -71971 -1686 -71970
rect -2298 -72098 -2171 -72082
rect -2298 -72222 -2194 -72098
rect -2298 -72238 -2171 -72222
rect -2727 -72350 -2405 -72349
rect -2727 -76480 -2726 -72350
rect -2406 -76480 -2405 -72350
rect -2727 -76481 -2405 -76480
rect -2618 -76859 -2514 -76481
rect -2298 -76592 -2251 -72238
rect -2187 -76592 -2171 -72238
rect -1899 -72349 -1795 -71971
rect -1579 -72082 -1532 -67728
rect -1468 -72082 -1452 -67728
rect -1180 -67839 -1076 -67461
rect -860 -67572 -813 -63218
rect -749 -67572 -733 -63218
rect -461 -63329 -357 -62951
rect -141 -63062 -94 -58708
rect -30 -63062 -14 -58708
rect 258 -58819 362 -58441
rect 578 -58552 625 -54198
rect 689 -58552 705 -54198
rect 977 -54309 1081 -53931
rect 1297 -54042 1344 -49688
rect 1408 -54042 1424 -49688
rect 1696 -49799 1800 -49421
rect 2016 -49532 2063 -45178
rect 2127 -49532 2143 -45178
rect 2415 -45289 2519 -44911
rect 2735 -45022 2782 -40668
rect 2846 -45022 2862 -40668
rect 2735 -45038 2862 -45022
rect 2735 -45162 2839 -45038
rect 2735 -45178 2862 -45162
rect 2306 -45290 2628 -45289
rect 2306 -49420 2307 -45290
rect 2627 -49420 2628 -45290
rect 2306 -49421 2628 -49420
rect 2016 -49548 2143 -49532
rect 2016 -49672 2120 -49548
rect 2016 -49688 2143 -49672
rect 1587 -49800 1909 -49799
rect 1587 -53930 1588 -49800
rect 1908 -53930 1909 -49800
rect 1587 -53931 1909 -53930
rect 1297 -54058 1424 -54042
rect 1297 -54182 1401 -54058
rect 1297 -54198 1424 -54182
rect 868 -54310 1190 -54309
rect 868 -58440 869 -54310
rect 1189 -58440 1190 -54310
rect 868 -58441 1190 -58440
rect 578 -58568 705 -58552
rect 578 -58692 682 -58568
rect 578 -58708 705 -58692
rect 149 -58820 471 -58819
rect 149 -62950 150 -58820
rect 470 -62950 471 -58820
rect 149 -62951 471 -62950
rect -141 -63078 -14 -63062
rect -141 -63202 -37 -63078
rect -141 -63218 -14 -63202
rect -570 -63330 -248 -63329
rect -570 -67460 -569 -63330
rect -249 -67460 -248 -63330
rect -570 -67461 -248 -67460
rect -860 -67588 -733 -67572
rect -860 -67712 -756 -67588
rect -860 -67728 -733 -67712
rect -1289 -67840 -967 -67839
rect -1289 -71970 -1288 -67840
rect -968 -71970 -967 -67840
rect -1289 -71971 -967 -71970
rect -1579 -72098 -1452 -72082
rect -1579 -72222 -1475 -72098
rect -1579 -72238 -1452 -72222
rect -2008 -72350 -1686 -72349
rect -2008 -76480 -2007 -72350
rect -1687 -76480 -1686 -72350
rect -2008 -76481 -1686 -76480
rect -2298 -76608 -2171 -76592
rect -2298 -76732 -2194 -76608
rect -2298 -76748 -2171 -76732
rect -2727 -76860 -2405 -76859
rect -2727 -80990 -2726 -76860
rect -2406 -80990 -2405 -76860
rect -2727 -80991 -2405 -80990
rect -2618 -81369 -2514 -80991
rect -2298 -81102 -2251 -76748
rect -2187 -81102 -2171 -76748
rect -1899 -76859 -1795 -76481
rect -1579 -76592 -1532 -72238
rect -1468 -76592 -1452 -72238
rect -1180 -72349 -1076 -71971
rect -860 -72082 -813 -67728
rect -749 -72082 -733 -67728
rect -461 -67839 -357 -67461
rect -141 -67572 -94 -63218
rect -30 -67572 -14 -63218
rect 258 -63329 362 -62951
rect 578 -63062 625 -58708
rect 689 -63062 705 -58708
rect 977 -58819 1081 -58441
rect 1297 -58552 1344 -54198
rect 1408 -58552 1424 -54198
rect 1696 -54309 1800 -53931
rect 2016 -54042 2063 -49688
rect 2127 -54042 2143 -49688
rect 2415 -49799 2519 -49421
rect 2735 -49532 2782 -45178
rect 2846 -49532 2862 -45178
rect 2735 -49548 2862 -49532
rect 2735 -49672 2839 -49548
rect 2735 -49688 2862 -49672
rect 2306 -49800 2628 -49799
rect 2306 -53930 2307 -49800
rect 2627 -53930 2628 -49800
rect 2306 -53931 2628 -53930
rect 2016 -54058 2143 -54042
rect 2016 -54182 2120 -54058
rect 2016 -54198 2143 -54182
rect 1587 -54310 1909 -54309
rect 1587 -58440 1588 -54310
rect 1908 -58440 1909 -54310
rect 1587 -58441 1909 -58440
rect 1297 -58568 1424 -58552
rect 1297 -58692 1401 -58568
rect 1297 -58708 1424 -58692
rect 868 -58820 1190 -58819
rect 868 -62950 869 -58820
rect 1189 -62950 1190 -58820
rect 868 -62951 1190 -62950
rect 578 -63078 705 -63062
rect 578 -63202 682 -63078
rect 578 -63218 705 -63202
rect 149 -63330 471 -63329
rect 149 -67460 150 -63330
rect 470 -67460 471 -63330
rect 149 -67461 471 -67460
rect -141 -67588 -14 -67572
rect -141 -67712 -37 -67588
rect -141 -67728 -14 -67712
rect -570 -67840 -248 -67839
rect -570 -71970 -569 -67840
rect -249 -71970 -248 -67840
rect -570 -71971 -248 -71970
rect -860 -72098 -733 -72082
rect -860 -72222 -756 -72098
rect -860 -72238 -733 -72222
rect -1289 -72350 -967 -72349
rect -1289 -76480 -1288 -72350
rect -968 -76480 -967 -72350
rect -1289 -76481 -967 -76480
rect -1579 -76608 -1452 -76592
rect -1579 -76732 -1475 -76608
rect -1579 -76748 -1452 -76732
rect -2008 -76860 -1686 -76859
rect -2008 -80990 -2007 -76860
rect -1687 -80990 -1686 -76860
rect -2008 -80991 -1686 -80990
rect -2298 -81118 -2171 -81102
rect -2298 -81242 -2194 -81118
rect -2298 -81258 -2171 -81242
rect -2727 -81370 -2405 -81369
rect -2727 -85500 -2726 -81370
rect -2406 -85500 -2405 -81370
rect -2727 -85501 -2405 -85500
rect -2618 -85879 -2514 -85501
rect -2298 -85612 -2251 -81258
rect -2187 -85612 -2171 -81258
rect -1899 -81369 -1795 -80991
rect -1579 -81102 -1532 -76748
rect -1468 -81102 -1452 -76748
rect -1180 -76859 -1076 -76481
rect -860 -76592 -813 -72238
rect -749 -76592 -733 -72238
rect -461 -72349 -357 -71971
rect -141 -72082 -94 -67728
rect -30 -72082 -14 -67728
rect 258 -67839 362 -67461
rect 578 -67572 625 -63218
rect 689 -67572 705 -63218
rect 977 -63329 1081 -62951
rect 1297 -63062 1344 -58708
rect 1408 -63062 1424 -58708
rect 1696 -58819 1800 -58441
rect 2016 -58552 2063 -54198
rect 2127 -58552 2143 -54198
rect 2415 -54309 2519 -53931
rect 2735 -54042 2782 -49688
rect 2846 -54042 2862 -49688
rect 2735 -54058 2862 -54042
rect 2735 -54182 2839 -54058
rect 2735 -54198 2862 -54182
rect 2306 -54310 2628 -54309
rect 2306 -58440 2307 -54310
rect 2627 -58440 2628 -54310
rect 2306 -58441 2628 -58440
rect 2016 -58568 2143 -58552
rect 2016 -58692 2120 -58568
rect 2016 -58708 2143 -58692
rect 1587 -58820 1909 -58819
rect 1587 -62950 1588 -58820
rect 1908 -62950 1909 -58820
rect 1587 -62951 1909 -62950
rect 1297 -63078 1424 -63062
rect 1297 -63202 1401 -63078
rect 1297 -63218 1424 -63202
rect 868 -63330 1190 -63329
rect 868 -67460 869 -63330
rect 1189 -67460 1190 -63330
rect 868 -67461 1190 -67460
rect 578 -67588 705 -67572
rect 578 -67712 682 -67588
rect 578 -67728 705 -67712
rect 149 -67840 471 -67839
rect 149 -71970 150 -67840
rect 470 -71970 471 -67840
rect 149 -71971 471 -71970
rect -141 -72098 -14 -72082
rect -141 -72222 -37 -72098
rect -141 -72238 -14 -72222
rect -570 -72350 -248 -72349
rect -570 -76480 -569 -72350
rect -249 -76480 -248 -72350
rect -570 -76481 -248 -76480
rect -860 -76608 -733 -76592
rect -860 -76732 -756 -76608
rect -860 -76748 -733 -76732
rect -1289 -76860 -967 -76859
rect -1289 -80990 -1288 -76860
rect -968 -80990 -967 -76860
rect -1289 -80991 -967 -80990
rect -1579 -81118 -1452 -81102
rect -1579 -81242 -1475 -81118
rect -1579 -81258 -1452 -81242
rect -2008 -81370 -1686 -81369
rect -2008 -85500 -2007 -81370
rect -1687 -85500 -1686 -81370
rect -2008 -85501 -1686 -85500
rect -2298 -85628 -2171 -85612
rect -2298 -85752 -2194 -85628
rect -2298 -85768 -2171 -85752
rect -2727 -85880 -2405 -85879
rect -2727 -90010 -2726 -85880
rect -2406 -90010 -2405 -85880
rect -2727 -90011 -2405 -90010
rect -2618 -90389 -2514 -90011
rect -2298 -90122 -2251 -85768
rect -2187 -90122 -2171 -85768
rect -1899 -85879 -1795 -85501
rect -1579 -85612 -1532 -81258
rect -1468 -85612 -1452 -81258
rect -1180 -81369 -1076 -80991
rect -860 -81102 -813 -76748
rect -749 -81102 -733 -76748
rect -461 -76859 -357 -76481
rect -141 -76592 -94 -72238
rect -30 -76592 -14 -72238
rect 258 -72349 362 -71971
rect 578 -72082 625 -67728
rect 689 -72082 705 -67728
rect 977 -67839 1081 -67461
rect 1297 -67572 1344 -63218
rect 1408 -67572 1424 -63218
rect 1696 -63329 1800 -62951
rect 2016 -63062 2063 -58708
rect 2127 -63062 2143 -58708
rect 2415 -58819 2519 -58441
rect 2735 -58552 2782 -54198
rect 2846 -58552 2862 -54198
rect 2735 -58568 2862 -58552
rect 2735 -58692 2839 -58568
rect 2735 -58708 2862 -58692
rect 2306 -58820 2628 -58819
rect 2306 -62950 2307 -58820
rect 2627 -62950 2628 -58820
rect 2306 -62951 2628 -62950
rect 2016 -63078 2143 -63062
rect 2016 -63202 2120 -63078
rect 2016 -63218 2143 -63202
rect 1587 -63330 1909 -63329
rect 1587 -67460 1588 -63330
rect 1908 -67460 1909 -63330
rect 1587 -67461 1909 -67460
rect 1297 -67588 1424 -67572
rect 1297 -67712 1401 -67588
rect 1297 -67728 1424 -67712
rect 868 -67840 1190 -67839
rect 868 -71970 869 -67840
rect 1189 -71970 1190 -67840
rect 868 -71971 1190 -71970
rect 578 -72098 705 -72082
rect 578 -72222 682 -72098
rect 578 -72238 705 -72222
rect 149 -72350 471 -72349
rect 149 -76480 150 -72350
rect 470 -76480 471 -72350
rect 149 -76481 471 -76480
rect -141 -76608 -14 -76592
rect -141 -76732 -37 -76608
rect -141 -76748 -14 -76732
rect -570 -76860 -248 -76859
rect -570 -80990 -569 -76860
rect -249 -80990 -248 -76860
rect -570 -80991 -248 -80990
rect -860 -81118 -733 -81102
rect -860 -81242 -756 -81118
rect -860 -81258 -733 -81242
rect -1289 -81370 -967 -81369
rect -1289 -85500 -1288 -81370
rect -968 -85500 -967 -81370
rect -1289 -85501 -967 -85500
rect -1579 -85628 -1452 -85612
rect -1579 -85752 -1475 -85628
rect -1579 -85768 -1452 -85752
rect -2008 -85880 -1686 -85879
rect -2008 -90010 -2007 -85880
rect -1687 -90010 -1686 -85880
rect -2008 -90011 -1686 -90010
rect -2298 -90138 -2171 -90122
rect -2298 -90262 -2194 -90138
rect -2298 -90278 -2171 -90262
rect -2727 -90390 -2405 -90389
rect -2727 -94520 -2726 -90390
rect -2406 -94520 -2405 -90390
rect -2727 -94521 -2405 -94520
rect -2618 -94899 -2514 -94521
rect -2298 -94632 -2251 -90278
rect -2187 -94632 -2171 -90278
rect -1899 -90389 -1795 -90011
rect -1579 -90122 -1532 -85768
rect -1468 -90122 -1452 -85768
rect -1180 -85879 -1076 -85501
rect -860 -85612 -813 -81258
rect -749 -85612 -733 -81258
rect -461 -81369 -357 -80991
rect -141 -81102 -94 -76748
rect -30 -81102 -14 -76748
rect 258 -76859 362 -76481
rect 578 -76592 625 -72238
rect 689 -76592 705 -72238
rect 977 -72349 1081 -71971
rect 1297 -72082 1344 -67728
rect 1408 -72082 1424 -67728
rect 1696 -67839 1800 -67461
rect 2016 -67572 2063 -63218
rect 2127 -67572 2143 -63218
rect 2415 -63329 2519 -62951
rect 2735 -63062 2782 -58708
rect 2846 -63062 2862 -58708
rect 2735 -63078 2862 -63062
rect 2735 -63202 2839 -63078
rect 2735 -63218 2862 -63202
rect 2306 -63330 2628 -63329
rect 2306 -67460 2307 -63330
rect 2627 -67460 2628 -63330
rect 2306 -67461 2628 -67460
rect 2016 -67588 2143 -67572
rect 2016 -67712 2120 -67588
rect 2016 -67728 2143 -67712
rect 1587 -67840 1909 -67839
rect 1587 -71970 1588 -67840
rect 1908 -71970 1909 -67840
rect 1587 -71971 1909 -71970
rect 1297 -72098 1424 -72082
rect 1297 -72222 1401 -72098
rect 1297 -72238 1424 -72222
rect 868 -72350 1190 -72349
rect 868 -76480 869 -72350
rect 1189 -76480 1190 -72350
rect 868 -76481 1190 -76480
rect 578 -76608 705 -76592
rect 578 -76732 682 -76608
rect 578 -76748 705 -76732
rect 149 -76860 471 -76859
rect 149 -80990 150 -76860
rect 470 -80990 471 -76860
rect 149 -80991 471 -80990
rect -141 -81118 -14 -81102
rect -141 -81242 -37 -81118
rect -141 -81258 -14 -81242
rect -570 -81370 -248 -81369
rect -570 -85500 -569 -81370
rect -249 -85500 -248 -81370
rect -570 -85501 -248 -85500
rect -860 -85628 -733 -85612
rect -860 -85752 -756 -85628
rect -860 -85768 -733 -85752
rect -1289 -85880 -967 -85879
rect -1289 -90010 -1288 -85880
rect -968 -90010 -967 -85880
rect -1289 -90011 -967 -90010
rect -1579 -90138 -1452 -90122
rect -1579 -90262 -1475 -90138
rect -1579 -90278 -1452 -90262
rect -2008 -90390 -1686 -90389
rect -2008 -94520 -2007 -90390
rect -1687 -94520 -1686 -90390
rect -2008 -94521 -1686 -94520
rect -2298 -94648 -2171 -94632
rect -2298 -94772 -2194 -94648
rect -2298 -94788 -2171 -94772
rect -2727 -94900 -2405 -94899
rect -2727 -99030 -2726 -94900
rect -2406 -99030 -2405 -94900
rect -2727 -99031 -2405 -99030
rect -2618 -99409 -2514 -99031
rect -2298 -99142 -2251 -94788
rect -2187 -99142 -2171 -94788
rect -1899 -94899 -1795 -94521
rect -1579 -94632 -1532 -90278
rect -1468 -94632 -1452 -90278
rect -1180 -90389 -1076 -90011
rect -860 -90122 -813 -85768
rect -749 -90122 -733 -85768
rect -461 -85879 -357 -85501
rect -141 -85612 -94 -81258
rect -30 -85612 -14 -81258
rect 258 -81369 362 -80991
rect 578 -81102 625 -76748
rect 689 -81102 705 -76748
rect 977 -76859 1081 -76481
rect 1297 -76592 1344 -72238
rect 1408 -76592 1424 -72238
rect 1696 -72349 1800 -71971
rect 2016 -72082 2063 -67728
rect 2127 -72082 2143 -67728
rect 2415 -67839 2519 -67461
rect 2735 -67572 2782 -63218
rect 2846 -67572 2862 -63218
rect 2735 -67588 2862 -67572
rect 2735 -67712 2839 -67588
rect 2735 -67728 2862 -67712
rect 2306 -67840 2628 -67839
rect 2306 -71970 2307 -67840
rect 2627 -71970 2628 -67840
rect 2306 -71971 2628 -71970
rect 2016 -72098 2143 -72082
rect 2016 -72222 2120 -72098
rect 2016 -72238 2143 -72222
rect 1587 -72350 1909 -72349
rect 1587 -76480 1588 -72350
rect 1908 -76480 1909 -72350
rect 1587 -76481 1909 -76480
rect 1297 -76608 1424 -76592
rect 1297 -76732 1401 -76608
rect 1297 -76748 1424 -76732
rect 868 -76860 1190 -76859
rect 868 -80990 869 -76860
rect 1189 -80990 1190 -76860
rect 868 -80991 1190 -80990
rect 578 -81118 705 -81102
rect 578 -81242 682 -81118
rect 578 -81258 705 -81242
rect 149 -81370 471 -81369
rect 149 -85500 150 -81370
rect 470 -85500 471 -81370
rect 149 -85501 471 -85500
rect -141 -85628 -14 -85612
rect -141 -85752 -37 -85628
rect -141 -85768 -14 -85752
rect -570 -85880 -248 -85879
rect -570 -90010 -569 -85880
rect -249 -90010 -248 -85880
rect -570 -90011 -248 -90010
rect -860 -90138 -733 -90122
rect -860 -90262 -756 -90138
rect -860 -90278 -733 -90262
rect -1289 -90390 -967 -90389
rect -1289 -94520 -1288 -90390
rect -968 -94520 -967 -90390
rect -1289 -94521 -967 -94520
rect -1579 -94648 -1452 -94632
rect -1579 -94772 -1475 -94648
rect -1579 -94788 -1452 -94772
rect -2008 -94900 -1686 -94899
rect -2008 -99030 -2007 -94900
rect -1687 -99030 -1686 -94900
rect -2008 -99031 -1686 -99030
rect -2298 -99158 -2171 -99142
rect -2298 -99282 -2194 -99158
rect -2298 -99298 -2171 -99282
rect -2727 -99410 -2405 -99409
rect -2727 -103540 -2726 -99410
rect -2406 -103540 -2405 -99410
rect -2727 -103541 -2405 -103540
rect -2618 -103919 -2514 -103541
rect -2298 -103652 -2251 -99298
rect -2187 -103652 -2171 -99298
rect -1899 -99409 -1795 -99031
rect -1579 -99142 -1532 -94788
rect -1468 -99142 -1452 -94788
rect -1180 -94899 -1076 -94521
rect -860 -94632 -813 -90278
rect -749 -94632 -733 -90278
rect -461 -90389 -357 -90011
rect -141 -90122 -94 -85768
rect -30 -90122 -14 -85768
rect 258 -85879 362 -85501
rect 578 -85612 625 -81258
rect 689 -85612 705 -81258
rect 977 -81369 1081 -80991
rect 1297 -81102 1344 -76748
rect 1408 -81102 1424 -76748
rect 1696 -76859 1800 -76481
rect 2016 -76592 2063 -72238
rect 2127 -76592 2143 -72238
rect 2415 -72349 2519 -71971
rect 2735 -72082 2782 -67728
rect 2846 -72082 2862 -67728
rect 2735 -72098 2862 -72082
rect 2735 -72222 2839 -72098
rect 2735 -72238 2862 -72222
rect 2306 -72350 2628 -72349
rect 2306 -76480 2307 -72350
rect 2627 -76480 2628 -72350
rect 2306 -76481 2628 -76480
rect 2016 -76608 2143 -76592
rect 2016 -76732 2120 -76608
rect 2016 -76748 2143 -76732
rect 1587 -76860 1909 -76859
rect 1587 -80990 1588 -76860
rect 1908 -80990 1909 -76860
rect 1587 -80991 1909 -80990
rect 1297 -81118 1424 -81102
rect 1297 -81242 1401 -81118
rect 1297 -81258 1424 -81242
rect 868 -81370 1190 -81369
rect 868 -85500 869 -81370
rect 1189 -85500 1190 -81370
rect 868 -85501 1190 -85500
rect 578 -85628 705 -85612
rect 578 -85752 682 -85628
rect 578 -85768 705 -85752
rect 149 -85880 471 -85879
rect 149 -90010 150 -85880
rect 470 -90010 471 -85880
rect 149 -90011 471 -90010
rect -141 -90138 -14 -90122
rect -141 -90262 -37 -90138
rect -141 -90278 -14 -90262
rect -570 -90390 -248 -90389
rect -570 -94520 -569 -90390
rect -249 -94520 -248 -90390
rect -570 -94521 -248 -94520
rect -860 -94648 -733 -94632
rect -860 -94772 -756 -94648
rect -860 -94788 -733 -94772
rect -1289 -94900 -967 -94899
rect -1289 -99030 -1288 -94900
rect -968 -99030 -967 -94900
rect -1289 -99031 -967 -99030
rect -1579 -99158 -1452 -99142
rect -1579 -99282 -1475 -99158
rect -1579 -99298 -1452 -99282
rect -2008 -99410 -1686 -99409
rect -2008 -103540 -2007 -99410
rect -1687 -103540 -1686 -99410
rect -2008 -103541 -1686 -103540
rect -2298 -103668 -2171 -103652
rect -2298 -103792 -2194 -103668
rect -2298 -103808 -2171 -103792
rect -2727 -103920 -2405 -103919
rect -2727 -108050 -2726 -103920
rect -2406 -108050 -2405 -103920
rect -2727 -108051 -2405 -108050
rect -2618 -108429 -2514 -108051
rect -2298 -108162 -2251 -103808
rect -2187 -108162 -2171 -103808
rect -1899 -103919 -1795 -103541
rect -1579 -103652 -1532 -99298
rect -1468 -103652 -1452 -99298
rect -1180 -99409 -1076 -99031
rect -860 -99142 -813 -94788
rect -749 -99142 -733 -94788
rect -461 -94899 -357 -94521
rect -141 -94632 -94 -90278
rect -30 -94632 -14 -90278
rect 258 -90389 362 -90011
rect 578 -90122 625 -85768
rect 689 -90122 705 -85768
rect 977 -85879 1081 -85501
rect 1297 -85612 1344 -81258
rect 1408 -85612 1424 -81258
rect 1696 -81369 1800 -80991
rect 2016 -81102 2063 -76748
rect 2127 -81102 2143 -76748
rect 2415 -76859 2519 -76481
rect 2735 -76592 2782 -72238
rect 2846 -76592 2862 -72238
rect 2735 -76608 2862 -76592
rect 2735 -76732 2839 -76608
rect 2735 -76748 2862 -76732
rect 2306 -76860 2628 -76859
rect 2306 -80990 2307 -76860
rect 2627 -80990 2628 -76860
rect 2306 -80991 2628 -80990
rect 2016 -81118 2143 -81102
rect 2016 -81242 2120 -81118
rect 2016 -81258 2143 -81242
rect 1587 -81370 1909 -81369
rect 1587 -85500 1588 -81370
rect 1908 -85500 1909 -81370
rect 1587 -85501 1909 -85500
rect 1297 -85628 1424 -85612
rect 1297 -85752 1401 -85628
rect 1297 -85768 1424 -85752
rect 868 -85880 1190 -85879
rect 868 -90010 869 -85880
rect 1189 -90010 1190 -85880
rect 868 -90011 1190 -90010
rect 578 -90138 705 -90122
rect 578 -90262 682 -90138
rect 578 -90278 705 -90262
rect 149 -90390 471 -90389
rect 149 -94520 150 -90390
rect 470 -94520 471 -90390
rect 149 -94521 471 -94520
rect -141 -94648 -14 -94632
rect -141 -94772 -37 -94648
rect -141 -94788 -14 -94772
rect -570 -94900 -248 -94899
rect -570 -99030 -569 -94900
rect -249 -99030 -248 -94900
rect -570 -99031 -248 -99030
rect -860 -99158 -733 -99142
rect -860 -99282 -756 -99158
rect -860 -99298 -733 -99282
rect -1289 -99410 -967 -99409
rect -1289 -103540 -1288 -99410
rect -968 -103540 -967 -99410
rect -1289 -103541 -967 -103540
rect -1579 -103668 -1452 -103652
rect -1579 -103792 -1475 -103668
rect -1579 -103808 -1452 -103792
rect -2008 -103920 -1686 -103919
rect -2008 -108050 -2007 -103920
rect -1687 -108050 -1686 -103920
rect -2008 -108051 -1686 -108050
rect -2298 -108178 -2171 -108162
rect -2298 -108302 -2194 -108178
rect -2298 -108318 -2171 -108302
rect -2727 -108430 -2405 -108429
rect -2727 -112560 -2726 -108430
rect -2406 -112560 -2405 -108430
rect -2727 -112561 -2405 -112560
rect -2618 -112939 -2514 -112561
rect -2298 -112672 -2251 -108318
rect -2187 -112672 -2171 -108318
rect -1899 -108429 -1795 -108051
rect -1579 -108162 -1532 -103808
rect -1468 -108162 -1452 -103808
rect -1180 -103919 -1076 -103541
rect -860 -103652 -813 -99298
rect -749 -103652 -733 -99298
rect -461 -99409 -357 -99031
rect -141 -99142 -94 -94788
rect -30 -99142 -14 -94788
rect 258 -94899 362 -94521
rect 578 -94632 625 -90278
rect 689 -94632 705 -90278
rect 977 -90389 1081 -90011
rect 1297 -90122 1344 -85768
rect 1408 -90122 1424 -85768
rect 1696 -85879 1800 -85501
rect 2016 -85612 2063 -81258
rect 2127 -85612 2143 -81258
rect 2415 -81369 2519 -80991
rect 2735 -81102 2782 -76748
rect 2846 -81102 2862 -76748
rect 2735 -81118 2862 -81102
rect 2735 -81242 2839 -81118
rect 2735 -81258 2862 -81242
rect 2306 -81370 2628 -81369
rect 2306 -85500 2307 -81370
rect 2627 -85500 2628 -81370
rect 2306 -85501 2628 -85500
rect 2016 -85628 2143 -85612
rect 2016 -85752 2120 -85628
rect 2016 -85768 2143 -85752
rect 1587 -85880 1909 -85879
rect 1587 -90010 1588 -85880
rect 1908 -90010 1909 -85880
rect 1587 -90011 1909 -90010
rect 1297 -90138 1424 -90122
rect 1297 -90262 1401 -90138
rect 1297 -90278 1424 -90262
rect 868 -90390 1190 -90389
rect 868 -94520 869 -90390
rect 1189 -94520 1190 -90390
rect 868 -94521 1190 -94520
rect 578 -94648 705 -94632
rect 578 -94772 682 -94648
rect 578 -94788 705 -94772
rect 149 -94900 471 -94899
rect 149 -99030 150 -94900
rect 470 -99030 471 -94900
rect 149 -99031 471 -99030
rect -141 -99158 -14 -99142
rect -141 -99282 -37 -99158
rect -141 -99298 -14 -99282
rect -570 -99410 -248 -99409
rect -570 -103540 -569 -99410
rect -249 -103540 -248 -99410
rect -570 -103541 -248 -103540
rect -860 -103668 -733 -103652
rect -860 -103792 -756 -103668
rect -860 -103808 -733 -103792
rect -1289 -103920 -967 -103919
rect -1289 -108050 -1288 -103920
rect -968 -108050 -967 -103920
rect -1289 -108051 -967 -108050
rect -1579 -108178 -1452 -108162
rect -1579 -108302 -1475 -108178
rect -1579 -108318 -1452 -108302
rect -2008 -108430 -1686 -108429
rect -2008 -112560 -2007 -108430
rect -1687 -112560 -1686 -108430
rect -2008 -112561 -1686 -112560
rect -2298 -112688 -2171 -112672
rect -2298 -112812 -2194 -112688
rect -2298 -112828 -2171 -112812
rect -2727 -112940 -2405 -112939
rect -2727 -117070 -2726 -112940
rect -2406 -117070 -2405 -112940
rect -2727 -117071 -2405 -117070
rect -2618 -117449 -2514 -117071
rect -2298 -117182 -2251 -112828
rect -2187 -117182 -2171 -112828
rect -1899 -112939 -1795 -112561
rect -1579 -112672 -1532 -108318
rect -1468 -112672 -1452 -108318
rect -1180 -108429 -1076 -108051
rect -860 -108162 -813 -103808
rect -749 -108162 -733 -103808
rect -461 -103919 -357 -103541
rect -141 -103652 -94 -99298
rect -30 -103652 -14 -99298
rect 258 -99409 362 -99031
rect 578 -99142 625 -94788
rect 689 -99142 705 -94788
rect 977 -94899 1081 -94521
rect 1297 -94632 1344 -90278
rect 1408 -94632 1424 -90278
rect 1696 -90389 1800 -90011
rect 2016 -90122 2063 -85768
rect 2127 -90122 2143 -85768
rect 2415 -85879 2519 -85501
rect 2735 -85612 2782 -81258
rect 2846 -85612 2862 -81258
rect 2735 -85628 2862 -85612
rect 2735 -85752 2839 -85628
rect 2735 -85768 2862 -85752
rect 2306 -85880 2628 -85879
rect 2306 -90010 2307 -85880
rect 2627 -90010 2628 -85880
rect 2306 -90011 2628 -90010
rect 2016 -90138 2143 -90122
rect 2016 -90262 2120 -90138
rect 2016 -90278 2143 -90262
rect 1587 -90390 1909 -90389
rect 1587 -94520 1588 -90390
rect 1908 -94520 1909 -90390
rect 1587 -94521 1909 -94520
rect 1297 -94648 1424 -94632
rect 1297 -94772 1401 -94648
rect 1297 -94788 1424 -94772
rect 868 -94900 1190 -94899
rect 868 -99030 869 -94900
rect 1189 -99030 1190 -94900
rect 868 -99031 1190 -99030
rect 578 -99158 705 -99142
rect 578 -99282 682 -99158
rect 578 -99298 705 -99282
rect 149 -99410 471 -99409
rect 149 -103540 150 -99410
rect 470 -103540 471 -99410
rect 149 -103541 471 -103540
rect -141 -103668 -14 -103652
rect -141 -103792 -37 -103668
rect -141 -103808 -14 -103792
rect -570 -103920 -248 -103919
rect -570 -108050 -569 -103920
rect -249 -108050 -248 -103920
rect -570 -108051 -248 -108050
rect -860 -108178 -733 -108162
rect -860 -108302 -756 -108178
rect -860 -108318 -733 -108302
rect -1289 -108430 -967 -108429
rect -1289 -112560 -1288 -108430
rect -968 -112560 -967 -108430
rect -1289 -112561 -967 -112560
rect -1579 -112688 -1452 -112672
rect -1579 -112812 -1475 -112688
rect -1579 -112828 -1452 -112812
rect -2008 -112940 -1686 -112939
rect -2008 -117070 -2007 -112940
rect -1687 -117070 -1686 -112940
rect -2008 -117071 -1686 -117070
rect -2298 -117198 -2171 -117182
rect -2298 -117322 -2194 -117198
rect -2298 -117338 -2171 -117322
rect -2727 -117450 -2405 -117449
rect -2727 -121580 -2726 -117450
rect -2406 -121580 -2405 -117450
rect -2727 -121581 -2405 -121580
rect -2618 -121959 -2514 -121581
rect -2298 -121692 -2251 -117338
rect -2187 -121692 -2171 -117338
rect -1899 -117449 -1795 -117071
rect -1579 -117182 -1532 -112828
rect -1468 -117182 -1452 -112828
rect -1180 -112939 -1076 -112561
rect -860 -112672 -813 -108318
rect -749 -112672 -733 -108318
rect -461 -108429 -357 -108051
rect -141 -108162 -94 -103808
rect -30 -108162 -14 -103808
rect 258 -103919 362 -103541
rect 578 -103652 625 -99298
rect 689 -103652 705 -99298
rect 977 -99409 1081 -99031
rect 1297 -99142 1344 -94788
rect 1408 -99142 1424 -94788
rect 1696 -94899 1800 -94521
rect 2016 -94632 2063 -90278
rect 2127 -94632 2143 -90278
rect 2415 -90389 2519 -90011
rect 2735 -90122 2782 -85768
rect 2846 -90122 2862 -85768
rect 2735 -90138 2862 -90122
rect 2735 -90262 2839 -90138
rect 2735 -90278 2862 -90262
rect 2306 -90390 2628 -90389
rect 2306 -94520 2307 -90390
rect 2627 -94520 2628 -90390
rect 2306 -94521 2628 -94520
rect 2016 -94648 2143 -94632
rect 2016 -94772 2120 -94648
rect 2016 -94788 2143 -94772
rect 1587 -94900 1909 -94899
rect 1587 -99030 1588 -94900
rect 1908 -99030 1909 -94900
rect 1587 -99031 1909 -99030
rect 1297 -99158 1424 -99142
rect 1297 -99282 1401 -99158
rect 1297 -99298 1424 -99282
rect 868 -99410 1190 -99409
rect 868 -103540 869 -99410
rect 1189 -103540 1190 -99410
rect 868 -103541 1190 -103540
rect 578 -103668 705 -103652
rect 578 -103792 682 -103668
rect 578 -103808 705 -103792
rect 149 -103920 471 -103919
rect 149 -108050 150 -103920
rect 470 -108050 471 -103920
rect 149 -108051 471 -108050
rect -141 -108178 -14 -108162
rect -141 -108302 -37 -108178
rect -141 -108318 -14 -108302
rect -570 -108430 -248 -108429
rect -570 -112560 -569 -108430
rect -249 -112560 -248 -108430
rect -570 -112561 -248 -112560
rect -860 -112688 -733 -112672
rect -860 -112812 -756 -112688
rect -860 -112828 -733 -112812
rect -1289 -112940 -967 -112939
rect -1289 -117070 -1288 -112940
rect -968 -117070 -967 -112940
rect -1289 -117071 -967 -117070
rect -1579 -117198 -1452 -117182
rect -1579 -117322 -1475 -117198
rect -1579 -117338 -1452 -117322
rect -2008 -117450 -1686 -117449
rect -2008 -121580 -2007 -117450
rect -1687 -121580 -1686 -117450
rect -2008 -121581 -1686 -121580
rect -2298 -121708 -2171 -121692
rect -2298 -121832 -2194 -121708
rect -2298 -121848 -2171 -121832
rect -2727 -121960 -2405 -121959
rect -2727 -126090 -2726 -121960
rect -2406 -126090 -2405 -121960
rect -2727 -126091 -2405 -126090
rect -2618 -126469 -2514 -126091
rect -2298 -126202 -2251 -121848
rect -2187 -126202 -2171 -121848
rect -1899 -121959 -1795 -121581
rect -1579 -121692 -1532 -117338
rect -1468 -121692 -1452 -117338
rect -1180 -117449 -1076 -117071
rect -860 -117182 -813 -112828
rect -749 -117182 -733 -112828
rect -461 -112939 -357 -112561
rect -141 -112672 -94 -108318
rect -30 -112672 -14 -108318
rect 258 -108429 362 -108051
rect 578 -108162 625 -103808
rect 689 -108162 705 -103808
rect 977 -103919 1081 -103541
rect 1297 -103652 1344 -99298
rect 1408 -103652 1424 -99298
rect 1696 -99409 1800 -99031
rect 2016 -99142 2063 -94788
rect 2127 -99142 2143 -94788
rect 2415 -94899 2519 -94521
rect 2735 -94632 2782 -90278
rect 2846 -94632 2862 -90278
rect 2735 -94648 2862 -94632
rect 2735 -94772 2839 -94648
rect 2735 -94788 2862 -94772
rect 2306 -94900 2628 -94899
rect 2306 -99030 2307 -94900
rect 2627 -99030 2628 -94900
rect 2306 -99031 2628 -99030
rect 2016 -99158 2143 -99142
rect 2016 -99282 2120 -99158
rect 2016 -99298 2143 -99282
rect 1587 -99410 1909 -99409
rect 1587 -103540 1588 -99410
rect 1908 -103540 1909 -99410
rect 1587 -103541 1909 -103540
rect 1297 -103668 1424 -103652
rect 1297 -103792 1401 -103668
rect 1297 -103808 1424 -103792
rect 868 -103920 1190 -103919
rect 868 -108050 869 -103920
rect 1189 -108050 1190 -103920
rect 868 -108051 1190 -108050
rect 578 -108178 705 -108162
rect 578 -108302 682 -108178
rect 578 -108318 705 -108302
rect 149 -108430 471 -108429
rect 149 -112560 150 -108430
rect 470 -112560 471 -108430
rect 149 -112561 471 -112560
rect -141 -112688 -14 -112672
rect -141 -112812 -37 -112688
rect -141 -112828 -14 -112812
rect -570 -112940 -248 -112939
rect -570 -117070 -569 -112940
rect -249 -117070 -248 -112940
rect -570 -117071 -248 -117070
rect -860 -117198 -733 -117182
rect -860 -117322 -756 -117198
rect -860 -117338 -733 -117322
rect -1289 -117450 -967 -117449
rect -1289 -121580 -1288 -117450
rect -968 -121580 -967 -117450
rect -1289 -121581 -967 -121580
rect -1579 -121708 -1452 -121692
rect -1579 -121832 -1475 -121708
rect -1579 -121848 -1452 -121832
rect -2008 -121960 -1686 -121959
rect -2008 -126090 -2007 -121960
rect -1687 -126090 -1686 -121960
rect -2008 -126091 -1686 -126090
rect -2298 -126218 -2171 -126202
rect -2298 -126342 -2194 -126218
rect -2298 -126358 -2171 -126342
rect -2727 -126470 -2405 -126469
rect -2727 -130600 -2726 -126470
rect -2406 -130600 -2405 -126470
rect -2727 -130601 -2405 -130600
rect -2618 -130979 -2514 -130601
rect -2298 -130712 -2251 -126358
rect -2187 -130712 -2171 -126358
rect -1899 -126469 -1795 -126091
rect -1579 -126202 -1532 -121848
rect -1468 -126202 -1452 -121848
rect -1180 -121959 -1076 -121581
rect -860 -121692 -813 -117338
rect -749 -121692 -733 -117338
rect -461 -117449 -357 -117071
rect -141 -117182 -94 -112828
rect -30 -117182 -14 -112828
rect 258 -112939 362 -112561
rect 578 -112672 625 -108318
rect 689 -112672 705 -108318
rect 977 -108429 1081 -108051
rect 1297 -108162 1344 -103808
rect 1408 -108162 1424 -103808
rect 1696 -103919 1800 -103541
rect 2016 -103652 2063 -99298
rect 2127 -103652 2143 -99298
rect 2415 -99409 2519 -99031
rect 2735 -99142 2782 -94788
rect 2846 -99142 2862 -94788
rect 2735 -99158 2862 -99142
rect 2735 -99282 2839 -99158
rect 2735 -99298 2862 -99282
rect 2306 -99410 2628 -99409
rect 2306 -103540 2307 -99410
rect 2627 -103540 2628 -99410
rect 2306 -103541 2628 -103540
rect 2016 -103668 2143 -103652
rect 2016 -103792 2120 -103668
rect 2016 -103808 2143 -103792
rect 1587 -103920 1909 -103919
rect 1587 -108050 1588 -103920
rect 1908 -108050 1909 -103920
rect 1587 -108051 1909 -108050
rect 1297 -108178 1424 -108162
rect 1297 -108302 1401 -108178
rect 1297 -108318 1424 -108302
rect 868 -108430 1190 -108429
rect 868 -112560 869 -108430
rect 1189 -112560 1190 -108430
rect 868 -112561 1190 -112560
rect 578 -112688 705 -112672
rect 578 -112812 682 -112688
rect 578 -112828 705 -112812
rect 149 -112940 471 -112939
rect 149 -117070 150 -112940
rect 470 -117070 471 -112940
rect 149 -117071 471 -117070
rect -141 -117198 -14 -117182
rect -141 -117322 -37 -117198
rect -141 -117338 -14 -117322
rect -570 -117450 -248 -117449
rect -570 -121580 -569 -117450
rect -249 -121580 -248 -117450
rect -570 -121581 -248 -121580
rect -860 -121708 -733 -121692
rect -860 -121832 -756 -121708
rect -860 -121848 -733 -121832
rect -1289 -121960 -967 -121959
rect -1289 -126090 -1288 -121960
rect -968 -126090 -967 -121960
rect -1289 -126091 -967 -126090
rect -1579 -126218 -1452 -126202
rect -1579 -126342 -1475 -126218
rect -1579 -126358 -1452 -126342
rect -2008 -126470 -1686 -126469
rect -2008 -130600 -2007 -126470
rect -1687 -130600 -1686 -126470
rect -2008 -130601 -1686 -130600
rect -2298 -130728 -2171 -130712
rect -2298 -130852 -2194 -130728
rect -2298 -130868 -2171 -130852
rect -2727 -130980 -2405 -130979
rect -2727 -135110 -2726 -130980
rect -2406 -135110 -2405 -130980
rect -2727 -135111 -2405 -135110
rect -2618 -135489 -2514 -135111
rect -2298 -135222 -2251 -130868
rect -2187 -135222 -2171 -130868
rect -1899 -130979 -1795 -130601
rect -1579 -130712 -1532 -126358
rect -1468 -130712 -1452 -126358
rect -1180 -126469 -1076 -126091
rect -860 -126202 -813 -121848
rect -749 -126202 -733 -121848
rect -461 -121959 -357 -121581
rect -141 -121692 -94 -117338
rect -30 -121692 -14 -117338
rect 258 -117449 362 -117071
rect 578 -117182 625 -112828
rect 689 -117182 705 -112828
rect 977 -112939 1081 -112561
rect 1297 -112672 1344 -108318
rect 1408 -112672 1424 -108318
rect 1696 -108429 1800 -108051
rect 2016 -108162 2063 -103808
rect 2127 -108162 2143 -103808
rect 2415 -103919 2519 -103541
rect 2735 -103652 2782 -99298
rect 2846 -103652 2862 -99298
rect 2735 -103668 2862 -103652
rect 2735 -103792 2839 -103668
rect 2735 -103808 2862 -103792
rect 2306 -103920 2628 -103919
rect 2306 -108050 2307 -103920
rect 2627 -108050 2628 -103920
rect 2306 -108051 2628 -108050
rect 2016 -108178 2143 -108162
rect 2016 -108302 2120 -108178
rect 2016 -108318 2143 -108302
rect 1587 -108430 1909 -108429
rect 1587 -112560 1588 -108430
rect 1908 -112560 1909 -108430
rect 1587 -112561 1909 -112560
rect 1297 -112688 1424 -112672
rect 1297 -112812 1401 -112688
rect 1297 -112828 1424 -112812
rect 868 -112940 1190 -112939
rect 868 -117070 869 -112940
rect 1189 -117070 1190 -112940
rect 868 -117071 1190 -117070
rect 578 -117198 705 -117182
rect 578 -117322 682 -117198
rect 578 -117338 705 -117322
rect 149 -117450 471 -117449
rect 149 -121580 150 -117450
rect 470 -121580 471 -117450
rect 149 -121581 471 -121580
rect -141 -121708 -14 -121692
rect -141 -121832 -37 -121708
rect -141 -121848 -14 -121832
rect -570 -121960 -248 -121959
rect -570 -126090 -569 -121960
rect -249 -126090 -248 -121960
rect -570 -126091 -248 -126090
rect -860 -126218 -733 -126202
rect -860 -126342 -756 -126218
rect -860 -126358 -733 -126342
rect -1289 -126470 -967 -126469
rect -1289 -130600 -1288 -126470
rect -968 -130600 -967 -126470
rect -1289 -130601 -967 -130600
rect -1579 -130728 -1452 -130712
rect -1579 -130852 -1475 -130728
rect -1579 -130868 -1452 -130852
rect -2008 -130980 -1686 -130979
rect -2008 -135110 -2007 -130980
rect -1687 -135110 -1686 -130980
rect -2008 -135111 -1686 -135110
rect -2298 -135238 -2171 -135222
rect -2298 -135362 -2194 -135238
rect -2298 -135378 -2171 -135362
rect -2727 -135490 -2405 -135489
rect -2727 -139620 -2726 -135490
rect -2406 -139620 -2405 -135490
rect -2727 -139621 -2405 -139620
rect -2618 -139999 -2514 -139621
rect -2298 -139732 -2251 -135378
rect -2187 -139732 -2171 -135378
rect -1899 -135489 -1795 -135111
rect -1579 -135222 -1532 -130868
rect -1468 -135222 -1452 -130868
rect -1180 -130979 -1076 -130601
rect -860 -130712 -813 -126358
rect -749 -130712 -733 -126358
rect -461 -126469 -357 -126091
rect -141 -126202 -94 -121848
rect -30 -126202 -14 -121848
rect 258 -121959 362 -121581
rect 578 -121692 625 -117338
rect 689 -121692 705 -117338
rect 977 -117449 1081 -117071
rect 1297 -117182 1344 -112828
rect 1408 -117182 1424 -112828
rect 1696 -112939 1800 -112561
rect 2016 -112672 2063 -108318
rect 2127 -112672 2143 -108318
rect 2415 -108429 2519 -108051
rect 2735 -108162 2782 -103808
rect 2846 -108162 2862 -103808
rect 2735 -108178 2862 -108162
rect 2735 -108302 2839 -108178
rect 2735 -108318 2862 -108302
rect 2306 -108430 2628 -108429
rect 2306 -112560 2307 -108430
rect 2627 -112560 2628 -108430
rect 2306 -112561 2628 -112560
rect 2016 -112688 2143 -112672
rect 2016 -112812 2120 -112688
rect 2016 -112828 2143 -112812
rect 1587 -112940 1909 -112939
rect 1587 -117070 1588 -112940
rect 1908 -117070 1909 -112940
rect 1587 -117071 1909 -117070
rect 1297 -117198 1424 -117182
rect 1297 -117322 1401 -117198
rect 1297 -117338 1424 -117322
rect 868 -117450 1190 -117449
rect 868 -121580 869 -117450
rect 1189 -121580 1190 -117450
rect 868 -121581 1190 -121580
rect 578 -121708 705 -121692
rect 578 -121832 682 -121708
rect 578 -121848 705 -121832
rect 149 -121960 471 -121959
rect 149 -126090 150 -121960
rect 470 -126090 471 -121960
rect 149 -126091 471 -126090
rect -141 -126218 -14 -126202
rect -141 -126342 -37 -126218
rect -141 -126358 -14 -126342
rect -570 -126470 -248 -126469
rect -570 -130600 -569 -126470
rect -249 -130600 -248 -126470
rect -570 -130601 -248 -130600
rect -860 -130728 -733 -130712
rect -860 -130852 -756 -130728
rect -860 -130868 -733 -130852
rect -1289 -130980 -967 -130979
rect -1289 -135110 -1288 -130980
rect -968 -135110 -967 -130980
rect -1289 -135111 -967 -135110
rect -1579 -135238 -1452 -135222
rect -1579 -135362 -1475 -135238
rect -1579 -135378 -1452 -135362
rect -2008 -135490 -1686 -135489
rect -2008 -139620 -2007 -135490
rect -1687 -139620 -1686 -135490
rect -2008 -139621 -1686 -139620
rect -2298 -139748 -2171 -139732
rect -2298 -139872 -2194 -139748
rect -2298 -139888 -2171 -139872
rect -2727 -140000 -2405 -139999
rect -2727 -144130 -2726 -140000
rect -2406 -144130 -2405 -140000
rect -2727 -144131 -2405 -144130
rect -2618 -144320 -2514 -144131
rect -2298 -144242 -2251 -139888
rect -2187 -144242 -2171 -139888
rect -1899 -139999 -1795 -139621
rect -1579 -139732 -1532 -135378
rect -1468 -139732 -1452 -135378
rect -1180 -135489 -1076 -135111
rect -860 -135222 -813 -130868
rect -749 -135222 -733 -130868
rect -461 -130979 -357 -130601
rect -141 -130712 -94 -126358
rect -30 -130712 -14 -126358
rect 258 -126469 362 -126091
rect 578 -126202 625 -121848
rect 689 -126202 705 -121848
rect 977 -121959 1081 -121581
rect 1297 -121692 1344 -117338
rect 1408 -121692 1424 -117338
rect 1696 -117449 1800 -117071
rect 2016 -117182 2063 -112828
rect 2127 -117182 2143 -112828
rect 2415 -112939 2519 -112561
rect 2735 -112672 2782 -108318
rect 2846 -112672 2862 -108318
rect 2735 -112688 2862 -112672
rect 2735 -112812 2839 -112688
rect 2735 -112828 2862 -112812
rect 2306 -112940 2628 -112939
rect 2306 -117070 2307 -112940
rect 2627 -117070 2628 -112940
rect 2306 -117071 2628 -117070
rect 2016 -117198 2143 -117182
rect 2016 -117322 2120 -117198
rect 2016 -117338 2143 -117322
rect 1587 -117450 1909 -117449
rect 1587 -121580 1588 -117450
rect 1908 -121580 1909 -117450
rect 1587 -121581 1909 -121580
rect 1297 -121708 1424 -121692
rect 1297 -121832 1401 -121708
rect 1297 -121848 1424 -121832
rect 868 -121960 1190 -121959
rect 868 -126090 869 -121960
rect 1189 -126090 1190 -121960
rect 868 -126091 1190 -126090
rect 578 -126218 705 -126202
rect 578 -126342 682 -126218
rect 578 -126358 705 -126342
rect 149 -126470 471 -126469
rect 149 -130600 150 -126470
rect 470 -130600 471 -126470
rect 149 -130601 471 -130600
rect -141 -130728 -14 -130712
rect -141 -130852 -37 -130728
rect -141 -130868 -14 -130852
rect -570 -130980 -248 -130979
rect -570 -135110 -569 -130980
rect -249 -135110 -248 -130980
rect -570 -135111 -248 -135110
rect -860 -135238 -733 -135222
rect -860 -135362 -756 -135238
rect -860 -135378 -733 -135362
rect -1289 -135490 -967 -135489
rect -1289 -139620 -1288 -135490
rect -968 -139620 -967 -135490
rect -1289 -139621 -967 -139620
rect -1579 -139748 -1452 -139732
rect -1579 -139872 -1475 -139748
rect -1579 -139888 -1452 -139872
rect -2008 -140000 -1686 -139999
rect -2008 -144130 -2007 -140000
rect -1687 -144130 -1686 -140000
rect -2008 -144131 -1686 -144130
rect -2298 -144258 -2171 -144242
rect -2298 -144320 -2194 -144258
rect -1899 -144320 -1795 -144131
rect -1579 -144242 -1532 -139888
rect -1468 -144242 -1452 -139888
rect -1180 -139999 -1076 -139621
rect -860 -139732 -813 -135378
rect -749 -139732 -733 -135378
rect -461 -135489 -357 -135111
rect -141 -135222 -94 -130868
rect -30 -135222 -14 -130868
rect 258 -130979 362 -130601
rect 578 -130712 625 -126358
rect 689 -130712 705 -126358
rect 977 -126469 1081 -126091
rect 1297 -126202 1344 -121848
rect 1408 -126202 1424 -121848
rect 1696 -121959 1800 -121581
rect 2016 -121692 2063 -117338
rect 2127 -121692 2143 -117338
rect 2415 -117449 2519 -117071
rect 2735 -117182 2782 -112828
rect 2846 -117182 2862 -112828
rect 2735 -117198 2862 -117182
rect 2735 -117322 2839 -117198
rect 2735 -117338 2862 -117322
rect 2306 -117450 2628 -117449
rect 2306 -121580 2307 -117450
rect 2627 -121580 2628 -117450
rect 2306 -121581 2628 -121580
rect 2016 -121708 2143 -121692
rect 2016 -121832 2120 -121708
rect 2016 -121848 2143 -121832
rect 1587 -121960 1909 -121959
rect 1587 -126090 1588 -121960
rect 1908 -126090 1909 -121960
rect 1587 -126091 1909 -126090
rect 1297 -126218 1424 -126202
rect 1297 -126342 1401 -126218
rect 1297 -126358 1424 -126342
rect 868 -126470 1190 -126469
rect 868 -130600 869 -126470
rect 1189 -130600 1190 -126470
rect 868 -130601 1190 -130600
rect 578 -130728 705 -130712
rect 578 -130852 682 -130728
rect 578 -130868 705 -130852
rect 149 -130980 471 -130979
rect 149 -135110 150 -130980
rect 470 -135110 471 -130980
rect 149 -135111 471 -135110
rect -141 -135238 -14 -135222
rect -141 -135362 -37 -135238
rect -141 -135378 -14 -135362
rect -570 -135490 -248 -135489
rect -570 -139620 -569 -135490
rect -249 -139620 -248 -135490
rect -570 -139621 -248 -139620
rect -860 -139748 -733 -139732
rect -860 -139872 -756 -139748
rect -860 -139888 -733 -139872
rect -1289 -140000 -967 -139999
rect -1289 -144130 -1288 -140000
rect -968 -144130 -967 -140000
rect -1289 -144131 -967 -144130
rect -1579 -144258 -1452 -144242
rect -1579 -144320 -1475 -144258
rect -1180 -144320 -1076 -144131
rect -860 -144242 -813 -139888
rect -749 -144242 -733 -139888
rect -461 -139999 -357 -139621
rect -141 -139732 -94 -135378
rect -30 -139732 -14 -135378
rect 258 -135489 362 -135111
rect 578 -135222 625 -130868
rect 689 -135222 705 -130868
rect 977 -130979 1081 -130601
rect 1297 -130712 1344 -126358
rect 1408 -130712 1424 -126358
rect 1696 -126469 1800 -126091
rect 2016 -126202 2063 -121848
rect 2127 -126202 2143 -121848
rect 2415 -121959 2519 -121581
rect 2735 -121692 2782 -117338
rect 2846 -121692 2862 -117338
rect 2735 -121708 2862 -121692
rect 2735 -121832 2839 -121708
rect 2735 -121848 2862 -121832
rect 2306 -121960 2628 -121959
rect 2306 -126090 2307 -121960
rect 2627 -126090 2628 -121960
rect 2306 -126091 2628 -126090
rect 2016 -126218 2143 -126202
rect 2016 -126342 2120 -126218
rect 2016 -126358 2143 -126342
rect 1587 -126470 1909 -126469
rect 1587 -130600 1588 -126470
rect 1908 -130600 1909 -126470
rect 1587 -130601 1909 -130600
rect 1297 -130728 1424 -130712
rect 1297 -130852 1401 -130728
rect 1297 -130868 1424 -130852
rect 868 -130980 1190 -130979
rect 868 -135110 869 -130980
rect 1189 -135110 1190 -130980
rect 868 -135111 1190 -135110
rect 578 -135238 705 -135222
rect 578 -135362 682 -135238
rect 578 -135378 705 -135362
rect 149 -135490 471 -135489
rect 149 -139620 150 -135490
rect 470 -139620 471 -135490
rect 149 -139621 471 -139620
rect -141 -139748 -14 -139732
rect -141 -139872 -37 -139748
rect -141 -139888 -14 -139872
rect -570 -140000 -248 -139999
rect -570 -144130 -569 -140000
rect -249 -144130 -248 -140000
rect -570 -144131 -248 -144130
rect -860 -144258 -733 -144242
rect -860 -144320 -756 -144258
rect -461 -144320 -357 -144131
rect -141 -144242 -94 -139888
rect -30 -144242 -14 -139888
rect 258 -139999 362 -139621
rect 578 -139732 625 -135378
rect 689 -139732 705 -135378
rect 977 -135489 1081 -135111
rect 1297 -135222 1344 -130868
rect 1408 -135222 1424 -130868
rect 1696 -130979 1800 -130601
rect 2016 -130712 2063 -126358
rect 2127 -130712 2143 -126358
rect 2415 -126469 2519 -126091
rect 2735 -126202 2782 -121848
rect 2846 -126202 2862 -121848
rect 2735 -126218 2862 -126202
rect 2735 -126342 2839 -126218
rect 2735 -126358 2862 -126342
rect 2306 -126470 2628 -126469
rect 2306 -130600 2307 -126470
rect 2627 -130600 2628 -126470
rect 2306 -130601 2628 -130600
rect 2016 -130728 2143 -130712
rect 2016 -130852 2120 -130728
rect 2016 -130868 2143 -130852
rect 1587 -130980 1909 -130979
rect 1587 -135110 1588 -130980
rect 1908 -135110 1909 -130980
rect 1587 -135111 1909 -135110
rect 1297 -135238 1424 -135222
rect 1297 -135362 1401 -135238
rect 1297 -135378 1424 -135362
rect 868 -135490 1190 -135489
rect 868 -139620 869 -135490
rect 1189 -139620 1190 -135490
rect 868 -139621 1190 -139620
rect 578 -139748 705 -139732
rect 578 -139872 682 -139748
rect 578 -139888 705 -139872
rect 149 -140000 471 -139999
rect 149 -144130 150 -140000
rect 470 -144130 471 -140000
rect 149 -144131 471 -144130
rect -141 -144258 -14 -144242
rect -141 -144320 -37 -144258
rect 258 -144320 362 -144131
rect 578 -144242 625 -139888
rect 689 -144242 705 -139888
rect 977 -139999 1081 -139621
rect 1297 -139732 1344 -135378
rect 1408 -139732 1424 -135378
rect 1696 -135489 1800 -135111
rect 2016 -135222 2063 -130868
rect 2127 -135222 2143 -130868
rect 2415 -130979 2519 -130601
rect 2735 -130712 2782 -126358
rect 2846 -130712 2862 -126358
rect 2735 -130728 2862 -130712
rect 2735 -130852 2839 -130728
rect 2735 -130868 2862 -130852
rect 2306 -130980 2628 -130979
rect 2306 -135110 2307 -130980
rect 2627 -135110 2628 -130980
rect 2306 -135111 2628 -135110
rect 2016 -135238 2143 -135222
rect 2016 -135362 2120 -135238
rect 2016 -135378 2143 -135362
rect 1587 -135490 1909 -135489
rect 1587 -139620 1588 -135490
rect 1908 -139620 1909 -135490
rect 1587 -139621 1909 -139620
rect 1297 -139748 1424 -139732
rect 1297 -139872 1401 -139748
rect 1297 -139888 1424 -139872
rect 868 -140000 1190 -139999
rect 868 -144130 869 -140000
rect 1189 -144130 1190 -140000
rect 868 -144131 1190 -144130
rect 578 -144258 705 -144242
rect 578 -144320 682 -144258
rect 977 -144320 1081 -144131
rect 1297 -144242 1344 -139888
rect 1408 -144242 1424 -139888
rect 1696 -139999 1800 -139621
rect 2016 -139732 2063 -135378
rect 2127 -139732 2143 -135378
rect 2415 -135489 2519 -135111
rect 2735 -135222 2782 -130868
rect 2846 -135222 2862 -130868
rect 2735 -135238 2862 -135222
rect 2735 -135362 2839 -135238
rect 2735 -135378 2862 -135362
rect 2306 -135490 2628 -135489
rect 2306 -139620 2307 -135490
rect 2627 -139620 2628 -135490
rect 2306 -139621 2628 -139620
rect 2016 -139748 2143 -139732
rect 2016 -139872 2120 -139748
rect 2016 -139888 2143 -139872
rect 1587 -140000 1909 -139999
rect 1587 -144130 1588 -140000
rect 1908 -144130 1909 -140000
rect 1587 -144131 1909 -144130
rect 1297 -144258 1424 -144242
rect 1297 -144320 1401 -144258
rect 1696 -144320 1800 -144131
rect 2016 -144242 2063 -139888
rect 2127 -144242 2143 -139888
rect 2415 -139999 2519 -139621
rect 2735 -139732 2782 -135378
rect 2846 -139732 2862 -135378
rect 2735 -139748 2862 -139732
rect 2735 -139872 2839 -139748
rect 2735 -139888 2862 -139872
rect 2306 -140000 2628 -139999
rect 2306 -144130 2307 -140000
rect 2627 -144130 2628 -140000
rect 2306 -144131 2628 -144130
rect 2016 -144258 2143 -144242
rect 2016 -144320 2120 -144258
rect 2415 -144320 2519 -144131
rect 2735 -144242 2782 -139888
rect 2846 -144242 2862 -139888
rect 2735 -144258 2862 -144242
rect 2735 -144320 2839 -144258
<< properties >>
string FIXED_BBOX 2167 139860 2767 144270
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 8 ny 64 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
