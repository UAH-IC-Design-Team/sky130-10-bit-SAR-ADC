magic
tech sky130A
magscale 1 2
timestamp 1666052912
<< metal4 >>
rect -2047 959 -949 1000
rect -2047 481 -1205 959
rect -969 481 -949 959
rect -2047 440 -949 481
rect -549 959 549 1000
rect -549 481 293 959
rect 529 481 549 959
rect -549 440 549 481
rect 949 959 2047 1000
rect 949 481 1791 959
rect 2027 481 2047 959
rect 949 440 2047 481
rect -2047 239 -949 280
rect -2047 -239 -1205 239
rect -969 -239 -949 239
rect -2047 -280 -949 -239
rect -549 239 549 280
rect -549 -239 293 239
rect 529 -239 549 239
rect -549 -280 549 -239
rect 949 239 2047 280
rect 949 -239 1791 239
rect 2027 -239 2047 239
rect 949 -280 2047 -239
rect -2047 -481 -949 -440
rect -2047 -959 -1205 -481
rect -969 -959 -949 -481
rect -2047 -1000 -949 -959
rect -549 -481 549 -440
rect -549 -959 293 -481
rect 529 -959 549 -481
rect -549 -1000 549 -959
rect 949 -481 2047 -440
rect 949 -959 1791 -481
rect 2027 -959 2047 -481
rect 949 -1000 2047 -959
<< via4 >>
rect -1205 481 -969 959
rect 293 481 529 959
rect 1791 481 2027 959
rect -1205 -239 -969 239
rect 293 -239 529 239
rect 1791 -239 2027 239
rect -1205 -959 -969 -481
rect 293 -959 529 -481
rect 1791 -959 2027 -481
<< mimcap2 >>
rect -1967 880 -1567 920
rect -1967 560 -1927 880
rect -1607 560 -1567 880
rect -1967 520 -1567 560
rect -469 880 -69 920
rect -469 560 -429 880
rect -109 560 -69 880
rect -469 520 -69 560
rect 1029 880 1429 920
rect 1029 560 1069 880
rect 1389 560 1429 880
rect 1029 520 1429 560
rect -1967 160 -1567 200
rect -1967 -160 -1927 160
rect -1607 -160 -1567 160
rect -1967 -200 -1567 -160
rect -469 160 -69 200
rect -469 -160 -429 160
rect -109 -160 -69 160
rect -469 -200 -69 -160
rect 1029 160 1429 200
rect 1029 -160 1069 160
rect 1389 -160 1429 160
rect 1029 -200 1429 -160
rect -1967 -560 -1567 -520
rect -1967 -880 -1927 -560
rect -1607 -880 -1567 -560
rect -1967 -920 -1567 -880
rect -469 -560 -69 -520
rect -469 -880 -429 -560
rect -109 -880 -69 -560
rect -469 -920 -69 -880
rect 1029 -560 1429 -520
rect 1029 -880 1069 -560
rect 1389 -880 1429 -560
rect 1029 -920 1429 -880
<< mimcap2contact >>
rect -1927 560 -1607 880
rect -429 560 -109 880
rect 1069 560 1389 880
rect -1927 -160 -1607 160
rect -429 -160 -109 160
rect 1069 -160 1389 160
rect -1927 -880 -1607 -560
rect -429 -880 -109 -560
rect 1069 -880 1389 -560
<< metal5 >>
rect -1927 904 -1607 1080
rect -1247 959 -927 1080
rect -1951 880 -1583 904
rect -1951 560 -1927 880
rect -1607 560 -1583 880
rect -1951 536 -1583 560
rect -1927 184 -1607 536
rect -1247 481 -1205 959
rect -969 481 -927 959
rect -429 904 -109 1080
rect 251 959 571 1080
rect -453 880 -85 904
rect -453 560 -429 880
rect -109 560 -85 880
rect -453 536 -85 560
rect -1247 239 -927 481
rect -1951 160 -1583 184
rect -1951 -160 -1927 160
rect -1607 -160 -1583 160
rect -1951 -184 -1583 -160
rect -1927 -536 -1607 -184
rect -1247 -239 -1205 239
rect -969 -239 -927 239
rect -429 184 -109 536
rect 251 481 293 959
rect 529 481 571 959
rect 1069 904 1389 1080
rect 1749 959 2069 1080
rect 1045 880 1413 904
rect 1045 560 1069 880
rect 1389 560 1413 880
rect 1045 536 1413 560
rect 251 239 571 481
rect -453 160 -85 184
rect -453 -160 -429 160
rect -109 -160 -85 160
rect -453 -184 -85 -160
rect -1247 -481 -927 -239
rect -1951 -560 -1583 -536
rect -1951 -880 -1927 -560
rect -1607 -880 -1583 -560
rect -1951 -904 -1583 -880
rect -1927 -1080 -1607 -904
rect -1247 -959 -1205 -481
rect -969 -959 -927 -481
rect -429 -536 -109 -184
rect 251 -239 293 239
rect 529 -239 571 239
rect 1069 184 1389 536
rect 1749 481 1791 959
rect 2027 481 2069 959
rect 1749 239 2069 481
rect 1045 160 1413 184
rect 1045 -160 1069 160
rect 1389 -160 1413 160
rect 1045 -184 1413 -160
rect 251 -481 571 -239
rect -453 -560 -85 -536
rect -453 -880 -429 -560
rect -109 -880 -85 -560
rect -453 -904 -85 -880
rect -1247 -1080 -927 -959
rect -429 -1080 -109 -904
rect 251 -959 293 -481
rect 529 -959 571 -481
rect 1069 -536 1389 -184
rect 1749 -239 1791 239
rect 2027 -239 2069 239
rect 1749 -481 2069 -239
rect 1045 -560 1413 -536
rect 1045 -880 1069 -560
rect 1389 -880 1413 -560
rect 1045 -904 1413 -880
rect 251 -1080 571 -959
rect 1069 -1080 1389 -904
rect 1749 -959 1791 -481
rect 2027 -959 2069 -481
rect 1749 -1080 2069 -959
<< properties >>
string FIXED_BBOX 949 440 1509 1000
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
