magic
tech sky130A
magscale 1 2
timestamp 1666651368
<< nmos >>
rect -687 -455 -657 455
rect -591 -455 -561 455
rect -495 -455 -465 455
rect -399 -455 -369 455
rect -303 -455 -273 455
rect -207 -455 -177 455
rect -111 -455 -81 455
rect -15 -455 15 455
rect 81 -455 111 455
rect 177 -455 207 455
rect 273 -455 303 455
rect 369 -455 399 455
rect 465 -455 495 455
rect 561 -455 591 455
rect 657 -455 687 455
<< ndiff >>
rect -749 443 -687 455
rect -749 -443 -737 443
rect -703 -443 -687 443
rect -749 -455 -687 -443
rect -657 443 -591 455
rect -657 -443 -641 443
rect -607 -443 -591 443
rect -657 -455 -591 -443
rect -561 443 -495 455
rect -561 -443 -545 443
rect -511 -443 -495 443
rect -561 -455 -495 -443
rect -465 443 -399 455
rect -465 -443 -449 443
rect -415 -443 -399 443
rect -465 -455 -399 -443
rect -369 443 -303 455
rect -369 -443 -353 443
rect -319 -443 -303 443
rect -369 -455 -303 -443
rect -273 443 -207 455
rect -273 -443 -257 443
rect -223 -443 -207 443
rect -273 -455 -207 -443
rect -177 443 -111 455
rect -177 -443 -161 443
rect -127 -443 -111 443
rect -177 -455 -111 -443
rect -81 443 -15 455
rect -81 -443 -65 443
rect -31 -443 -15 443
rect -81 -455 -15 -443
rect 15 443 81 455
rect 15 -443 31 443
rect 65 -443 81 443
rect 15 -455 81 -443
rect 111 443 177 455
rect 111 -443 127 443
rect 161 -443 177 443
rect 111 -455 177 -443
rect 207 443 273 455
rect 207 -443 223 443
rect 257 -443 273 443
rect 207 -455 273 -443
rect 303 443 369 455
rect 303 -443 319 443
rect 353 -443 369 443
rect 303 -455 369 -443
rect 399 443 465 455
rect 399 -443 415 443
rect 449 -443 465 443
rect 399 -455 465 -443
rect 495 443 561 455
rect 495 -443 511 443
rect 545 -443 561 443
rect 495 -455 561 -443
rect 591 443 657 455
rect 591 -443 607 443
rect 641 -443 657 443
rect 591 -455 657 -443
rect 687 443 749 455
rect 687 -443 703 443
rect 737 -443 749 443
rect 687 -455 749 -443
<< ndiffc >>
rect -737 -443 -703 443
rect -641 -443 -607 443
rect -545 -443 -511 443
rect -449 -443 -415 443
rect -353 -443 -319 443
rect -257 -443 -223 443
rect -161 -443 -127 443
rect -65 -443 -31 443
rect 31 -443 65 443
rect 127 -443 161 443
rect 223 -443 257 443
rect 319 -443 353 443
rect 415 -443 449 443
rect 511 -443 545 443
rect 607 -443 641 443
rect 703 -443 737 443
<< poly >>
rect -687 455 -657 484
rect -591 455 -561 484
rect -495 455 -465 484
rect -399 455 -369 484
rect -303 455 -273 484
rect -207 455 -177 484
rect -111 455 -81 484
rect -15 455 15 484
rect 81 455 111 484
rect 177 455 207 484
rect 273 455 303 484
rect 369 455 399 484
rect 465 455 495 484
rect 561 455 591 484
rect 657 455 687 484
rect -687 -476 -657 -455
rect -591 -476 -561 -455
rect -495 -476 -465 -455
rect -399 -476 -369 -455
rect -303 -476 -273 -455
rect -207 -476 -177 -455
rect -111 -476 -81 -455
rect -15 -476 15 -455
rect 81 -476 111 -455
rect 177 -476 207 -455
rect 273 -476 303 -455
rect 369 -476 399 -455
rect 465 -476 495 -455
rect 561 -476 591 -455
rect 657 -476 687 -455
rect -708 -493 705 -476
rect -708 -527 -689 -493
rect -655 -527 -594 -493
rect -560 -527 -497 -493
rect -463 -527 -394 -493
rect -360 -527 -305 -493
rect -271 -527 -204 -493
rect -170 -527 -113 -493
rect -79 -527 -14 -493
rect 20 -527 79 -493
rect 113 -527 176 -493
rect 210 -527 271 -493
rect 305 -527 375 -493
rect 409 -527 463 -493
rect 497 -527 565 -493
rect 599 -527 655 -493
rect 689 -527 705 -493
rect -708 -543 705 -527
<< polycont >>
rect -689 -527 -655 -493
rect -594 -527 -560 -493
rect -497 -527 -463 -493
rect -394 -527 -360 -493
rect -305 -527 -271 -493
rect -204 -527 -170 -493
rect -113 -527 -79 -493
rect -14 -527 20 -493
rect 79 -527 113 -493
rect 176 -527 210 -493
rect 271 -527 305 -493
rect 375 -527 409 -493
rect 463 -527 497 -493
rect 565 -527 599 -493
rect 655 -527 689 -493
<< locali >>
rect -737 443 -703 459
rect -737 -459 -703 -443
rect -641 443 -607 459
rect -641 -459 -607 -443
rect -545 443 -511 459
rect -545 -459 -511 -443
rect -449 443 -415 459
rect -449 -459 -415 -443
rect -353 443 -319 459
rect -353 -459 -319 -443
rect -257 443 -223 459
rect -257 -459 -223 -443
rect -161 443 -127 459
rect -161 -459 -127 -443
rect -65 443 -31 459
rect -65 -459 -31 -443
rect 31 443 65 459
rect 31 -459 65 -443
rect 127 443 161 459
rect 127 -459 161 -443
rect 223 443 257 459
rect 223 -459 257 -443
rect 319 443 353 459
rect 319 -459 353 -443
rect 415 443 449 459
rect 415 -459 449 -443
rect 511 443 545 459
rect 511 -459 545 -443
rect 607 443 641 459
rect 607 -459 641 -443
rect 703 443 737 459
rect 703 -459 737 -443
rect -708 -527 -689 -493
rect -655 -527 -594 -493
rect -560 -527 -497 -493
rect -463 -527 -394 -493
rect -360 -527 -305 -493
rect -271 -527 -204 -493
rect -170 -527 -113 -493
rect -79 -527 -14 -493
rect 20 -527 79 -493
rect 113 -527 176 -493
rect 210 -527 271 -493
rect 305 -527 375 -493
rect 409 -527 463 -493
rect 497 -527 565 -493
rect 599 -527 655 -493
rect 689 -527 705 -493
<< viali >>
rect -737 -426 -703 -72
rect -641 72 -607 426
rect -545 -426 -511 -72
rect -449 72 -415 426
rect -353 -426 -319 -72
rect -257 72 -223 426
rect -161 -426 -127 -72
rect -65 72 -31 426
rect 31 -426 65 -72
rect 127 72 161 426
rect 223 -426 257 -72
rect 319 72 353 426
rect 415 -426 449 -72
rect 511 72 545 426
rect 607 -426 641 -72
rect 703 72 737 426
rect -689 -527 -655 -493
rect -594 -527 -560 -493
rect -497 -527 -463 -493
rect -394 -527 -360 -493
rect -305 -527 -271 -493
rect -204 -527 -170 -493
rect -113 -527 -79 -493
rect -14 -527 20 -493
rect 79 -527 113 -493
rect 176 -527 210 -493
rect 271 -527 305 -493
rect 375 -527 409 -493
rect 463 -527 497 -493
rect 565 -527 599 -493
rect 655 -527 689 -493
<< metal1 >>
rect -647 426 -601 438
rect -647 72 -641 426
rect -607 72 -601 426
rect -647 60 -601 72
rect -455 426 -409 438
rect -455 72 -449 426
rect -415 72 -409 426
rect -455 60 -409 72
rect -263 426 -217 438
rect -263 72 -257 426
rect -223 72 -217 426
rect -263 60 -217 72
rect -71 426 -25 438
rect -71 72 -65 426
rect -31 72 -25 426
rect -71 60 -25 72
rect 121 426 167 438
rect 121 72 127 426
rect 161 72 167 426
rect 121 60 167 72
rect 313 426 359 438
rect 313 72 319 426
rect 353 72 359 426
rect 313 60 359 72
rect 505 426 551 438
rect 505 72 511 426
rect 545 72 551 426
rect 505 60 551 72
rect 697 426 743 438
rect 697 72 703 426
rect 737 72 743 426
rect 697 60 743 72
rect -743 -72 -697 -60
rect -743 -426 -737 -72
rect -703 -426 -697 -72
rect -743 -438 -697 -426
rect -551 -72 -505 -60
rect -551 -426 -545 -72
rect -511 -426 -505 -72
rect -551 -438 -505 -426
rect -359 -72 -313 -60
rect -359 -426 -353 -72
rect -319 -426 -313 -72
rect -359 -438 -313 -426
rect -167 -72 -121 -60
rect -167 -426 -161 -72
rect -127 -426 -121 -72
rect -167 -438 -121 -426
rect 25 -72 71 -60
rect 25 -426 31 -72
rect 65 -426 71 -72
rect 25 -438 71 -426
rect 217 -72 263 -60
rect 217 -426 223 -72
rect 257 -426 263 -72
rect 217 -438 263 -426
rect 409 -72 455 -60
rect 409 -426 415 -72
rect 449 -426 455 -72
rect 409 -438 455 -426
rect 601 -72 647 -60
rect 601 -426 607 -72
rect 641 -426 647 -72
rect 601 -438 647 -426
rect -708 -493 701 -487
rect -708 -527 -689 -493
rect -655 -527 -594 -493
rect -560 -527 -497 -493
rect -463 -527 -394 -493
rect -360 -527 -305 -493
rect -271 -527 -204 -493
rect -170 -527 -113 -493
rect -79 -527 -14 -493
rect 20 -527 79 -493
rect 113 -527 176 -493
rect 210 -527 271 -493
rect 305 -527 375 -493
rect 409 -527 463 -493
rect 497 -527 565 -493
rect 599 -527 655 -493
rect 689 -527 701 -493
rect -708 -533 701 -527
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.55 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
