magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< error_p >>
rect -789 13580 -729 17990
rect -709 13580 -649 17990
rect -70 13580 -10 17990
rect 10 13580 70 17990
rect 649 13580 709 17990
rect 729 13580 789 17990
rect -789 9070 -729 13480
rect -709 9070 -649 13480
rect -70 9070 -10 13480
rect 10 9070 70 13480
rect 649 9070 709 13480
rect 729 9070 789 13480
rect -789 4560 -729 8970
rect -709 4560 -649 8970
rect -70 4560 -10 8970
rect 10 4560 70 8970
rect 649 4560 709 8970
rect 729 4560 789 8970
rect -789 50 -729 4460
rect -709 50 -649 4460
rect -70 50 -10 4460
rect 10 50 70 4460
rect 649 50 709 4460
rect 729 50 789 4460
rect -789 -4460 -729 -50
rect -709 -4460 -649 -50
rect -70 -4460 -10 -50
rect 10 -4460 70 -50
rect 649 -4460 709 -50
rect 729 -4460 789 -50
rect -789 -8970 -729 -4560
rect -709 -8970 -649 -4560
rect -70 -8970 -10 -4560
rect 10 -8970 70 -4560
rect 649 -8970 709 -4560
rect 729 -8970 789 -4560
rect -789 -13480 -729 -9070
rect -709 -13480 -649 -9070
rect -70 -13480 -10 -9070
rect 10 -13480 70 -9070
rect 649 -13480 709 -9070
rect 729 -13480 789 -9070
rect -789 -17990 -729 -13580
rect -709 -17990 -649 -13580
rect -70 -17990 -10 -13580
rect 10 -17990 70 -13580
rect 649 -17990 709 -13580
rect 729 -17990 789 -13580
<< metal3 >>
rect -1428 17962 -729 17990
rect -1428 13608 -813 17962
rect -749 13608 -729 17962
rect -1428 13580 -729 13608
rect -709 17962 -10 17990
rect -709 13608 -94 17962
rect -30 13608 -10 17962
rect -709 13580 -10 13608
rect 10 17962 709 17990
rect 10 13608 625 17962
rect 689 13608 709 17962
rect 10 13580 709 13608
rect 729 17962 1428 17990
rect 729 13608 1344 17962
rect 1408 13608 1428 17962
rect 729 13580 1428 13608
rect -1428 13452 -729 13480
rect -1428 9098 -813 13452
rect -749 9098 -729 13452
rect -1428 9070 -729 9098
rect -709 13452 -10 13480
rect -709 9098 -94 13452
rect -30 9098 -10 13452
rect -709 9070 -10 9098
rect 10 13452 709 13480
rect 10 9098 625 13452
rect 689 9098 709 13452
rect 10 9070 709 9098
rect 729 13452 1428 13480
rect 729 9098 1344 13452
rect 1408 9098 1428 13452
rect 729 9070 1428 9098
rect -1428 8942 -729 8970
rect -1428 4588 -813 8942
rect -749 4588 -729 8942
rect -1428 4560 -729 4588
rect -709 8942 -10 8970
rect -709 4588 -94 8942
rect -30 4588 -10 8942
rect -709 4560 -10 4588
rect 10 8942 709 8970
rect 10 4588 625 8942
rect 689 4588 709 8942
rect 10 4560 709 4588
rect 729 8942 1428 8970
rect 729 4588 1344 8942
rect 1408 4588 1428 8942
rect 729 4560 1428 4588
rect -1428 4432 -729 4460
rect -1428 78 -813 4432
rect -749 78 -729 4432
rect -1428 50 -729 78
rect -709 4432 -10 4460
rect -709 78 -94 4432
rect -30 78 -10 4432
rect -709 50 -10 78
rect 10 4432 709 4460
rect 10 78 625 4432
rect 689 78 709 4432
rect 10 50 709 78
rect 729 4432 1428 4460
rect 729 78 1344 4432
rect 1408 78 1428 4432
rect 729 50 1428 78
rect -1428 -78 -729 -50
rect -1428 -4432 -813 -78
rect -749 -4432 -729 -78
rect -1428 -4460 -729 -4432
rect -709 -78 -10 -50
rect -709 -4432 -94 -78
rect -30 -4432 -10 -78
rect -709 -4460 -10 -4432
rect 10 -78 709 -50
rect 10 -4432 625 -78
rect 689 -4432 709 -78
rect 10 -4460 709 -4432
rect 729 -78 1428 -50
rect 729 -4432 1344 -78
rect 1408 -4432 1428 -78
rect 729 -4460 1428 -4432
rect -1428 -4588 -729 -4560
rect -1428 -8942 -813 -4588
rect -749 -8942 -729 -4588
rect -1428 -8970 -729 -8942
rect -709 -4588 -10 -4560
rect -709 -8942 -94 -4588
rect -30 -8942 -10 -4588
rect -709 -8970 -10 -8942
rect 10 -4588 709 -4560
rect 10 -8942 625 -4588
rect 689 -8942 709 -4588
rect 10 -8970 709 -8942
rect 729 -4588 1428 -4560
rect 729 -8942 1344 -4588
rect 1408 -8942 1428 -4588
rect 729 -8970 1428 -8942
rect -1428 -9098 -729 -9070
rect -1428 -13452 -813 -9098
rect -749 -13452 -729 -9098
rect -1428 -13480 -729 -13452
rect -709 -9098 -10 -9070
rect -709 -13452 -94 -9098
rect -30 -13452 -10 -9098
rect -709 -13480 -10 -13452
rect 10 -9098 709 -9070
rect 10 -13452 625 -9098
rect 689 -13452 709 -9098
rect 10 -13480 709 -13452
rect 729 -9098 1428 -9070
rect 729 -13452 1344 -9098
rect 1408 -13452 1428 -9098
rect 729 -13480 1428 -13452
rect -1428 -13608 -729 -13580
rect -1428 -17962 -813 -13608
rect -749 -17962 -729 -13608
rect -1428 -17990 -729 -17962
rect -709 -13608 -10 -13580
rect -709 -17962 -94 -13608
rect -30 -17962 -10 -13608
rect -709 -17990 -10 -17962
rect 10 -13608 709 -13580
rect 10 -17962 625 -13608
rect 689 -17962 709 -13608
rect 10 -17990 709 -17962
rect 729 -13608 1428 -13580
rect 729 -17962 1344 -13608
rect 1408 -17962 1428 -13608
rect 729 -17990 1428 -17962
<< via3 >>
rect -813 13608 -749 17962
rect -94 13608 -30 17962
rect 625 13608 689 17962
rect 1344 13608 1408 17962
rect -813 9098 -749 13452
rect -94 9098 -30 13452
rect 625 9098 689 13452
rect 1344 9098 1408 13452
rect -813 4588 -749 8942
rect -94 4588 -30 8942
rect 625 4588 689 8942
rect 1344 4588 1408 8942
rect -813 78 -749 4432
rect -94 78 -30 4432
rect 625 78 689 4432
rect 1344 78 1408 4432
rect -813 -4432 -749 -78
rect -94 -4432 -30 -78
rect 625 -4432 689 -78
rect 1344 -4432 1408 -78
rect -813 -8942 -749 -4588
rect -94 -8942 -30 -4588
rect 625 -8942 689 -4588
rect 1344 -8942 1408 -4588
rect -813 -13452 -749 -9098
rect -94 -13452 -30 -9098
rect 625 -13452 689 -9098
rect 1344 -13452 1408 -9098
rect -813 -17962 -749 -13608
rect -94 -17962 -30 -13608
rect 625 -17962 689 -13608
rect 1344 -17962 1408 -13608
<< mimcap >>
rect -1328 17850 -928 17890
rect -1328 13720 -1288 17850
rect -968 13720 -928 17850
rect -1328 13680 -928 13720
rect -609 17850 -209 17890
rect -609 13720 -569 17850
rect -249 13720 -209 17850
rect -609 13680 -209 13720
rect 110 17850 510 17890
rect 110 13720 150 17850
rect 470 13720 510 17850
rect 110 13680 510 13720
rect 829 17850 1229 17890
rect 829 13720 869 17850
rect 1189 13720 1229 17850
rect 829 13680 1229 13720
rect -1328 13340 -928 13380
rect -1328 9210 -1288 13340
rect -968 9210 -928 13340
rect -1328 9170 -928 9210
rect -609 13340 -209 13380
rect -609 9210 -569 13340
rect -249 9210 -209 13340
rect -609 9170 -209 9210
rect 110 13340 510 13380
rect 110 9210 150 13340
rect 470 9210 510 13340
rect 110 9170 510 9210
rect 829 13340 1229 13380
rect 829 9210 869 13340
rect 1189 9210 1229 13340
rect 829 9170 1229 9210
rect -1328 8830 -928 8870
rect -1328 4700 -1288 8830
rect -968 4700 -928 8830
rect -1328 4660 -928 4700
rect -609 8830 -209 8870
rect -609 4700 -569 8830
rect -249 4700 -209 8830
rect -609 4660 -209 4700
rect 110 8830 510 8870
rect 110 4700 150 8830
rect 470 4700 510 8830
rect 110 4660 510 4700
rect 829 8830 1229 8870
rect 829 4700 869 8830
rect 1189 4700 1229 8830
rect 829 4660 1229 4700
rect -1328 4320 -928 4360
rect -1328 190 -1288 4320
rect -968 190 -928 4320
rect -1328 150 -928 190
rect -609 4320 -209 4360
rect -609 190 -569 4320
rect -249 190 -209 4320
rect -609 150 -209 190
rect 110 4320 510 4360
rect 110 190 150 4320
rect 470 190 510 4320
rect 110 150 510 190
rect 829 4320 1229 4360
rect 829 190 869 4320
rect 1189 190 1229 4320
rect 829 150 1229 190
rect -1328 -190 -928 -150
rect -1328 -4320 -1288 -190
rect -968 -4320 -928 -190
rect -1328 -4360 -928 -4320
rect -609 -190 -209 -150
rect -609 -4320 -569 -190
rect -249 -4320 -209 -190
rect -609 -4360 -209 -4320
rect 110 -190 510 -150
rect 110 -4320 150 -190
rect 470 -4320 510 -190
rect 110 -4360 510 -4320
rect 829 -190 1229 -150
rect 829 -4320 869 -190
rect 1189 -4320 1229 -190
rect 829 -4360 1229 -4320
rect -1328 -4700 -928 -4660
rect -1328 -8830 -1288 -4700
rect -968 -8830 -928 -4700
rect -1328 -8870 -928 -8830
rect -609 -4700 -209 -4660
rect -609 -8830 -569 -4700
rect -249 -8830 -209 -4700
rect -609 -8870 -209 -8830
rect 110 -4700 510 -4660
rect 110 -8830 150 -4700
rect 470 -8830 510 -4700
rect 110 -8870 510 -8830
rect 829 -4700 1229 -4660
rect 829 -8830 869 -4700
rect 1189 -8830 1229 -4700
rect 829 -8870 1229 -8830
rect -1328 -9210 -928 -9170
rect -1328 -13340 -1288 -9210
rect -968 -13340 -928 -9210
rect -1328 -13380 -928 -13340
rect -609 -9210 -209 -9170
rect -609 -13340 -569 -9210
rect -249 -13340 -209 -9210
rect -609 -13380 -209 -13340
rect 110 -9210 510 -9170
rect 110 -13340 150 -9210
rect 470 -13340 510 -9210
rect 110 -13380 510 -13340
rect 829 -9210 1229 -9170
rect 829 -13340 869 -9210
rect 1189 -13340 1229 -9210
rect 829 -13380 1229 -13340
rect -1328 -13720 -928 -13680
rect -1328 -17850 -1288 -13720
rect -968 -17850 -928 -13720
rect -1328 -17890 -928 -17850
rect -609 -13720 -209 -13680
rect -609 -17850 -569 -13720
rect -249 -17850 -209 -13720
rect -609 -17890 -209 -17850
rect 110 -13720 510 -13680
rect 110 -17850 150 -13720
rect 470 -17850 510 -13720
rect 110 -17890 510 -17850
rect 829 -13720 1229 -13680
rect 829 -17850 869 -13720
rect 1189 -17850 1229 -13720
rect 829 -17890 1229 -17850
<< mimcapcontact >>
rect -1288 13720 -968 17850
rect -569 13720 -249 17850
rect 150 13720 470 17850
rect 869 13720 1189 17850
rect -1288 9210 -968 13340
rect -569 9210 -249 13340
rect 150 9210 470 13340
rect 869 9210 1189 13340
rect -1288 4700 -968 8830
rect -569 4700 -249 8830
rect 150 4700 470 8830
rect 869 4700 1189 8830
rect -1288 190 -968 4320
rect -569 190 -249 4320
rect 150 190 470 4320
rect 869 190 1189 4320
rect -1288 -4320 -968 -190
rect -569 -4320 -249 -190
rect 150 -4320 470 -190
rect 869 -4320 1189 -190
rect -1288 -8830 -968 -4700
rect -569 -8830 -249 -4700
rect 150 -8830 470 -4700
rect 869 -8830 1189 -4700
rect -1288 -13340 -968 -9210
rect -569 -13340 -249 -9210
rect 150 -13340 470 -9210
rect 869 -13340 1189 -9210
rect -1288 -17850 -968 -13720
rect -569 -17850 -249 -13720
rect 150 -17850 470 -13720
rect 869 -17850 1189 -13720
<< metal4 >>
rect -1180 17851 -1076 18040
rect -860 17978 -756 18040
rect -860 17962 -733 17978
rect -1289 17850 -967 17851
rect -1289 13720 -1288 17850
rect -968 13720 -967 17850
rect -1289 13719 -967 13720
rect -1180 13341 -1076 13719
rect -860 13608 -813 17962
rect -749 13608 -733 17962
rect -461 17851 -357 18040
rect -141 17978 -37 18040
rect -141 17962 -14 17978
rect -570 17850 -248 17851
rect -570 13720 -569 17850
rect -249 13720 -248 17850
rect -570 13719 -248 13720
rect -860 13592 -733 13608
rect -860 13468 -756 13592
rect -860 13452 -733 13468
rect -1289 13340 -967 13341
rect -1289 9210 -1288 13340
rect -968 9210 -967 13340
rect -1289 9209 -967 9210
rect -1180 8831 -1076 9209
rect -860 9098 -813 13452
rect -749 9098 -733 13452
rect -461 13341 -357 13719
rect -141 13608 -94 17962
rect -30 13608 -14 17962
rect 258 17851 362 18040
rect 578 17978 682 18040
rect 578 17962 705 17978
rect 149 17850 471 17851
rect 149 13720 150 17850
rect 470 13720 471 17850
rect 149 13719 471 13720
rect -141 13592 -14 13608
rect -141 13468 -37 13592
rect -141 13452 -14 13468
rect -570 13340 -248 13341
rect -570 9210 -569 13340
rect -249 9210 -248 13340
rect -570 9209 -248 9210
rect -860 9082 -733 9098
rect -860 8958 -756 9082
rect -860 8942 -733 8958
rect -1289 8830 -967 8831
rect -1289 4700 -1288 8830
rect -968 4700 -967 8830
rect -1289 4699 -967 4700
rect -1180 4321 -1076 4699
rect -860 4588 -813 8942
rect -749 4588 -733 8942
rect -461 8831 -357 9209
rect -141 9098 -94 13452
rect -30 9098 -14 13452
rect 258 13341 362 13719
rect 578 13608 625 17962
rect 689 13608 705 17962
rect 977 17851 1081 18040
rect 1297 17978 1401 18040
rect 1297 17962 1424 17978
rect 868 17850 1190 17851
rect 868 13720 869 17850
rect 1189 13720 1190 17850
rect 868 13719 1190 13720
rect 578 13592 705 13608
rect 578 13468 682 13592
rect 578 13452 705 13468
rect 149 13340 471 13341
rect 149 9210 150 13340
rect 470 9210 471 13340
rect 149 9209 471 9210
rect -141 9082 -14 9098
rect -141 8958 -37 9082
rect -141 8942 -14 8958
rect -570 8830 -248 8831
rect -570 4700 -569 8830
rect -249 4700 -248 8830
rect -570 4699 -248 4700
rect -860 4572 -733 4588
rect -860 4448 -756 4572
rect -860 4432 -733 4448
rect -1289 4320 -967 4321
rect -1289 190 -1288 4320
rect -968 190 -967 4320
rect -1289 189 -967 190
rect -1180 -189 -1076 189
rect -860 78 -813 4432
rect -749 78 -733 4432
rect -461 4321 -357 4699
rect -141 4588 -94 8942
rect -30 4588 -14 8942
rect 258 8831 362 9209
rect 578 9098 625 13452
rect 689 9098 705 13452
rect 977 13341 1081 13719
rect 1297 13608 1344 17962
rect 1408 13608 1424 17962
rect 1297 13592 1424 13608
rect 1297 13468 1401 13592
rect 1297 13452 1424 13468
rect 868 13340 1190 13341
rect 868 9210 869 13340
rect 1189 9210 1190 13340
rect 868 9209 1190 9210
rect 578 9082 705 9098
rect 578 8958 682 9082
rect 578 8942 705 8958
rect 149 8830 471 8831
rect 149 4700 150 8830
rect 470 4700 471 8830
rect 149 4699 471 4700
rect -141 4572 -14 4588
rect -141 4448 -37 4572
rect -141 4432 -14 4448
rect -570 4320 -248 4321
rect -570 190 -569 4320
rect -249 190 -248 4320
rect -570 189 -248 190
rect -860 62 -733 78
rect -860 -62 -756 62
rect -860 -78 -733 -62
rect -1289 -190 -967 -189
rect -1289 -4320 -1288 -190
rect -968 -4320 -967 -190
rect -1289 -4321 -967 -4320
rect -1180 -4699 -1076 -4321
rect -860 -4432 -813 -78
rect -749 -4432 -733 -78
rect -461 -189 -357 189
rect -141 78 -94 4432
rect -30 78 -14 4432
rect 258 4321 362 4699
rect 578 4588 625 8942
rect 689 4588 705 8942
rect 977 8831 1081 9209
rect 1297 9098 1344 13452
rect 1408 9098 1424 13452
rect 1297 9082 1424 9098
rect 1297 8958 1401 9082
rect 1297 8942 1424 8958
rect 868 8830 1190 8831
rect 868 4700 869 8830
rect 1189 4700 1190 8830
rect 868 4699 1190 4700
rect 578 4572 705 4588
rect 578 4448 682 4572
rect 578 4432 705 4448
rect 149 4320 471 4321
rect 149 190 150 4320
rect 470 190 471 4320
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -4320 -569 -190
rect -249 -4320 -248 -190
rect -570 -4321 -248 -4320
rect -860 -4448 -733 -4432
rect -860 -4572 -756 -4448
rect -860 -4588 -733 -4572
rect -1289 -4700 -967 -4699
rect -1289 -8830 -1288 -4700
rect -968 -8830 -967 -4700
rect -1289 -8831 -967 -8830
rect -1180 -9209 -1076 -8831
rect -860 -8942 -813 -4588
rect -749 -8942 -733 -4588
rect -461 -4699 -357 -4321
rect -141 -4432 -94 -78
rect -30 -4432 -14 -78
rect 258 -189 362 189
rect 578 78 625 4432
rect 689 78 705 4432
rect 977 4321 1081 4699
rect 1297 4588 1344 8942
rect 1408 4588 1424 8942
rect 1297 4572 1424 4588
rect 1297 4448 1401 4572
rect 1297 4432 1424 4448
rect 868 4320 1190 4321
rect 868 190 869 4320
rect 1189 190 1190 4320
rect 868 189 1190 190
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -4320 150 -190
rect 470 -4320 471 -190
rect 149 -4321 471 -4320
rect -141 -4448 -14 -4432
rect -141 -4572 -37 -4448
rect -141 -4588 -14 -4572
rect -570 -4700 -248 -4699
rect -570 -8830 -569 -4700
rect -249 -8830 -248 -4700
rect -570 -8831 -248 -8830
rect -860 -8958 -733 -8942
rect -860 -9082 -756 -8958
rect -860 -9098 -733 -9082
rect -1289 -9210 -967 -9209
rect -1289 -13340 -1288 -9210
rect -968 -13340 -967 -9210
rect -1289 -13341 -967 -13340
rect -1180 -13719 -1076 -13341
rect -860 -13452 -813 -9098
rect -749 -13452 -733 -9098
rect -461 -9209 -357 -8831
rect -141 -8942 -94 -4588
rect -30 -8942 -14 -4588
rect 258 -4699 362 -4321
rect 578 -4432 625 -78
rect 689 -4432 705 -78
rect 977 -189 1081 189
rect 1297 78 1344 4432
rect 1408 78 1424 4432
rect 1297 62 1424 78
rect 1297 -62 1401 62
rect 1297 -78 1424 -62
rect 868 -190 1190 -189
rect 868 -4320 869 -190
rect 1189 -4320 1190 -190
rect 868 -4321 1190 -4320
rect 578 -4448 705 -4432
rect 578 -4572 682 -4448
rect 578 -4588 705 -4572
rect 149 -4700 471 -4699
rect 149 -8830 150 -4700
rect 470 -8830 471 -4700
rect 149 -8831 471 -8830
rect -141 -8958 -14 -8942
rect -141 -9082 -37 -8958
rect -141 -9098 -14 -9082
rect -570 -9210 -248 -9209
rect -570 -13340 -569 -9210
rect -249 -13340 -248 -9210
rect -570 -13341 -248 -13340
rect -860 -13468 -733 -13452
rect -860 -13592 -756 -13468
rect -860 -13608 -733 -13592
rect -1289 -13720 -967 -13719
rect -1289 -17850 -1288 -13720
rect -968 -17850 -967 -13720
rect -1289 -17851 -967 -17850
rect -1180 -18040 -1076 -17851
rect -860 -17962 -813 -13608
rect -749 -17962 -733 -13608
rect -461 -13719 -357 -13341
rect -141 -13452 -94 -9098
rect -30 -13452 -14 -9098
rect 258 -9209 362 -8831
rect 578 -8942 625 -4588
rect 689 -8942 705 -4588
rect 977 -4699 1081 -4321
rect 1297 -4432 1344 -78
rect 1408 -4432 1424 -78
rect 1297 -4448 1424 -4432
rect 1297 -4572 1401 -4448
rect 1297 -4588 1424 -4572
rect 868 -4700 1190 -4699
rect 868 -8830 869 -4700
rect 1189 -8830 1190 -4700
rect 868 -8831 1190 -8830
rect 578 -8958 705 -8942
rect 578 -9082 682 -8958
rect 578 -9098 705 -9082
rect 149 -9210 471 -9209
rect 149 -13340 150 -9210
rect 470 -13340 471 -9210
rect 149 -13341 471 -13340
rect -141 -13468 -14 -13452
rect -141 -13592 -37 -13468
rect -141 -13608 -14 -13592
rect -570 -13720 -248 -13719
rect -570 -17850 -569 -13720
rect -249 -17850 -248 -13720
rect -570 -17851 -248 -17850
rect -860 -17978 -733 -17962
rect -860 -18040 -756 -17978
rect -461 -18040 -357 -17851
rect -141 -17962 -94 -13608
rect -30 -17962 -14 -13608
rect 258 -13719 362 -13341
rect 578 -13452 625 -9098
rect 689 -13452 705 -9098
rect 977 -9209 1081 -8831
rect 1297 -8942 1344 -4588
rect 1408 -8942 1424 -4588
rect 1297 -8958 1424 -8942
rect 1297 -9082 1401 -8958
rect 1297 -9098 1424 -9082
rect 868 -9210 1190 -9209
rect 868 -13340 869 -9210
rect 1189 -13340 1190 -9210
rect 868 -13341 1190 -13340
rect 578 -13468 705 -13452
rect 578 -13592 682 -13468
rect 578 -13608 705 -13592
rect 149 -13720 471 -13719
rect 149 -17850 150 -13720
rect 470 -17850 471 -13720
rect 149 -17851 471 -17850
rect -141 -17978 -14 -17962
rect -141 -18040 -37 -17978
rect 258 -18040 362 -17851
rect 578 -17962 625 -13608
rect 689 -17962 705 -13608
rect 977 -13719 1081 -13341
rect 1297 -13452 1344 -9098
rect 1408 -13452 1424 -9098
rect 1297 -13468 1424 -13452
rect 1297 -13592 1401 -13468
rect 1297 -13608 1424 -13592
rect 868 -13720 1190 -13719
rect 868 -17850 869 -13720
rect 1189 -17850 1190 -13720
rect 868 -17851 1190 -17850
rect 578 -17978 705 -17962
rect 578 -18040 682 -17978
rect 977 -18040 1081 -17851
rect 1297 -17962 1344 -13608
rect 1408 -17962 1424 -13608
rect 1297 -17978 1424 -17962
rect 1297 -18040 1401 -17978
<< properties >>
string FIXED_BBOX 729 13580 1329 17990
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
