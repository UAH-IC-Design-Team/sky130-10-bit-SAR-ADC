magic
tech sky130A
magscale 1 2
timestamp 1666486738
<< error_p >>
rect -29 1095 29 1101
rect -29 1061 -17 1095
rect -29 1055 29 1061
rect -29 637 29 643
rect -29 603 -17 637
rect -29 597 29 603
rect -29 529 29 535
rect -29 495 -17 529
rect -29 489 29 495
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -495 29 -489
rect -29 -529 -17 -495
rect -29 -535 29 -529
rect -29 -603 29 -597
rect -29 -637 -17 -603
rect -29 -643 29 -637
rect -29 -1061 29 -1055
rect -29 -1095 -17 -1061
rect -29 -1101 29 -1095
<< nwell >>
rect -211 -1233 211 1233
<< pmos >>
rect -15 684 15 1014
rect -15 118 15 448
rect -15 -448 15 -118
rect -15 -1014 15 -684
<< pdiff >>
rect -73 1002 -15 1014
rect -73 696 -61 1002
rect -27 696 -15 1002
rect -73 684 -15 696
rect 15 1002 73 1014
rect 15 696 27 1002
rect 61 696 73 1002
rect 15 684 73 696
rect -73 436 -15 448
rect -73 130 -61 436
rect -27 130 -15 436
rect -73 118 -15 130
rect 15 436 73 448
rect 15 130 27 436
rect 61 130 73 436
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -436 -61 -130
rect -27 -436 -15 -130
rect -73 -448 -15 -436
rect 15 -130 73 -118
rect 15 -436 27 -130
rect 61 -436 73 -130
rect 15 -448 73 -436
rect -73 -696 -15 -684
rect -73 -1002 -61 -696
rect -27 -1002 -15 -696
rect -73 -1014 -15 -1002
rect 15 -696 73 -684
rect 15 -1002 27 -696
rect 61 -1002 73 -696
rect 15 -1014 73 -1002
<< pdiffc >>
rect -61 696 -27 1002
rect 27 696 61 1002
rect -61 130 -27 436
rect 27 130 61 436
rect -61 -436 -27 -130
rect 27 -436 61 -130
rect -61 -1002 -27 -696
rect 27 -1002 61 -696
<< nsubdiff >>
rect -175 1163 -79 1197
rect 79 1163 175 1197
rect -175 1101 -141 1163
rect 141 1101 175 1163
rect -175 -1163 -141 -1101
rect 141 -1163 175 -1101
rect -175 -1197 -79 -1163
rect 79 -1197 175 -1163
<< nsubdiffcont >>
rect -79 1163 79 1197
rect -175 -1101 -141 1101
rect 141 -1101 175 1101
rect -79 -1197 79 -1163
<< poly >>
rect -33 1095 33 1111
rect -33 1061 -17 1095
rect 17 1061 33 1095
rect -33 1045 33 1061
rect -15 1014 15 1045
rect -15 653 15 684
rect -33 637 33 653
rect -33 603 -17 637
rect 17 603 33 637
rect -33 587 33 603
rect -33 529 33 545
rect -33 495 -17 529
rect 17 495 33 529
rect -33 479 33 495
rect -15 448 15 479
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -479 15 -448
rect -33 -495 33 -479
rect -33 -529 -17 -495
rect 17 -529 33 -495
rect -33 -545 33 -529
rect -33 -603 33 -587
rect -33 -637 -17 -603
rect 17 -637 33 -603
rect -33 -653 33 -637
rect -15 -684 15 -653
rect -15 -1045 15 -1014
rect -33 -1061 33 -1045
rect -33 -1095 -17 -1061
rect 17 -1095 33 -1061
rect -33 -1111 33 -1095
<< polycont >>
rect -17 1061 17 1095
rect -17 603 17 637
rect -17 495 17 529
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -529 17 -495
rect -17 -637 17 -603
rect -17 -1095 17 -1061
<< locali >>
rect -175 1163 -79 1197
rect 79 1163 175 1197
rect -175 1101 -141 1163
rect 141 1101 175 1163
rect -33 1061 -17 1095
rect 17 1061 33 1095
rect -61 1002 -27 1018
rect -61 680 -27 696
rect 27 1002 61 1018
rect 27 680 61 696
rect -33 603 -17 637
rect 17 603 33 637
rect -33 495 -17 529
rect 17 495 33 529
rect -61 436 -27 452
rect -61 114 -27 130
rect 27 436 61 452
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -452 -27 -436
rect 27 -130 61 -114
rect 27 -452 61 -436
rect -33 -529 -17 -495
rect 17 -529 33 -495
rect -33 -637 -17 -603
rect 17 -637 33 -603
rect -61 -696 -27 -680
rect -61 -1018 -27 -1002
rect 27 -696 61 -680
rect 27 -1018 61 -1002
rect -33 -1095 -17 -1061
rect 17 -1095 33 -1061
rect -175 -1163 -141 -1101
rect 141 -1163 175 -1101
rect -175 -1197 -79 -1163
rect 79 -1197 175 -1163
<< viali >>
rect -17 1061 17 1095
rect -61 696 -27 1002
rect 27 696 61 1002
rect -17 603 17 637
rect -17 495 17 529
rect -61 130 -27 436
rect 27 130 61 436
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -436 -27 -130
rect 27 -436 61 -130
rect -17 -529 17 -495
rect -17 -637 17 -603
rect -61 -1002 -27 -696
rect 27 -1002 61 -696
rect -17 -1095 17 -1061
<< metal1 >>
rect -29 1095 29 1101
rect -29 1061 -17 1095
rect 17 1061 29 1095
rect -29 1055 29 1061
rect -67 1002 -21 1014
rect -67 696 -61 1002
rect -27 696 -21 1002
rect -67 684 -21 696
rect 21 1002 67 1014
rect 21 696 27 1002
rect 61 696 67 1002
rect 21 684 67 696
rect -29 637 29 643
rect -29 603 -17 637
rect 17 603 29 637
rect -29 597 29 603
rect -29 529 29 535
rect -29 495 -17 529
rect 17 495 29 529
rect -29 489 29 495
rect -67 436 -21 448
rect -67 130 -61 436
rect -27 130 -21 436
rect -67 118 -21 130
rect 21 436 67 448
rect 21 130 27 436
rect 61 130 67 436
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -436 -61 -130
rect -27 -436 -21 -130
rect -67 -448 -21 -436
rect 21 -130 67 -118
rect 21 -436 27 -130
rect 61 -436 67 -130
rect 21 -448 67 -436
rect -29 -495 29 -489
rect -29 -529 -17 -495
rect 17 -529 29 -495
rect -29 -535 29 -529
rect -29 -603 29 -597
rect -29 -637 -17 -603
rect 17 -637 29 -603
rect -29 -643 29 -637
rect -67 -696 -21 -684
rect -67 -1002 -61 -696
rect -27 -1002 -21 -696
rect -67 -1014 -21 -1002
rect 21 -696 67 -684
rect 21 -1002 27 -696
rect 61 -1002 67 -696
rect 21 -1014 67 -1002
rect -29 -1061 29 -1055
rect -29 -1095 -17 -1061
rect 17 -1095 29 -1061
rect -29 -1101 29 -1095
<< properties >>
string FIXED_BBOX -158 -1180 158 1180
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
