** CONTROLLER flat netlist
*.PININFO CLK:I SW_N_SP[9..1]:O VSS:B VDD:B RESET:I VCMP:I SW_N[8..1]:O SW_P_SP[9..1]:O SW_P[8..1]:O
*+ BIT[10..1]:O DONE:O SW_SAMPLE:O
*--------BEGIN_X95->SKY130_FD_SC_HD__OR4_2
X95 CYCLE1 CYCLE2 CYCLE3 CYCLE4 VSS VSS VDD VDD NET2  SKY130_FD_SC_HD__OR4_2
*--------END___X95->SKY130_FD_SC_HD__OR4_2
*--------BEGIN_X96->SKY130_FD_SC_HD__OR4_2
X96 CYCLE5 CYCLE6 CYCLE7 CYCLE8 VSS VSS VDD VDD NET3  SKY130_FD_SC_HD__OR4_2
*--------END___X96->SKY130_FD_SC_HD__OR4_2
*--------BEGIN_X97->SKY130_FD_SC_HD__OR4_2
X97 CYCLE9 CYCLE10 CYCLE11 CYCLE12 VSS VSS VDD VDD NET5  SKY130_FD_SC_HD__OR4_2
*--------END___X97->SKY130_FD_SC_HD__OR4_2
*--------BEGIN_X3->DEC
*.PININFO VDD:B BIT[10..1]:O VSS:B RESET_B:I DUMP_BUS:I DONE:O RAW_BIT[13..1]:I
*--------BEGIN_X3_X62->SKY130_FD_SC_HD__FA_1
X62_X3 RAW_BIT2 RAW_BIT1 X3_NET1 VSS VSS VDD VDD X3_NET16 X3_NET2  SKY130_FD_SC_HD__FA_1
*--------END___X3_X62->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X64->SKY130_FD_SC_HD__FA_1
X64_X3 RAW_BIT3 RAW_BIT1 X3_NET4 VSS VSS VDD VDD X3_NET1 X3_NET3  SKY130_FD_SC_HD__FA_1
*--------END___X3_X64->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X67->SKY130_FD_SC_HD__DFRTP_1
X67_X3 CYCLE31 X3_NET2 RESET VSS VSS VDD VDD BIT2  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X67->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X68->SKY130_FD_SC_HD__DFRTP_1
X68_X3 CYCLE31 X3_NET3 RESET VSS VSS VDD VDD BIT3  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X68->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X65->SKY130_FD_SC_HD__FA_1
X65_X3 RAW_BIT5 RAW_BIT4 X3_NET5 VSS VSS VDD VDD X3_NET4 X3_NET6  SKY130_FD_SC_HD__FA_1
*--------END___X3_X65->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X69->SKY130_FD_SC_HD__FA_1
X69_X3 RAW_BIT6 RAW_BIT4 X3_NET8 VSS VSS VDD VDD X3_NET5 X3_NET7  SKY130_FD_SC_HD__FA_1
*--------END___X3_X69->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X70->SKY130_FD_SC_HD__DFRTP_1
X70_X3 CYCLE31 X3_NET6 RESET VSS VSS VDD VDD BIT4  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X70->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X71->SKY130_FD_SC_HD__DFRTP_1
X71_X3 CYCLE31 X3_NET7 RESET VSS VSS VDD VDD BIT5  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X71->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X72->SKY130_FD_SC_HD__FA_1
X72_X3 RAW_BIT7 RAW_BIT4 X3_NET9 VSS VSS VDD VDD X3_NET8 X3_NET10  SKY130_FD_SC_HD__FA_1
*--------END___X3_X72->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X73->SKY130_FD_SC_HD__FA_1
X73_X3 RAW_BIT9 RAW_BIT8 X3_NET12 VSS VSS VDD VDD X3_NET9 X3_NET11  SKY130_FD_SC_HD__FA_1
*--------END___X3_X73->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X74->SKY130_FD_SC_HD__DFRTP_1
X74_X3 CYCLE31 X3_NET10 RESET VSS VSS VDD VDD BIT6  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X74->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X75->SKY130_FD_SC_HD__DFRTP_1
X75_X3 CYCLE31 X3_NET11 RESET VSS VSS VDD VDD BIT7  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X75->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X76->SKY130_FD_SC_HD__FA_1
X76_X3 RAW_BIT10 RAW_BIT8 X3_NET13 VSS VSS VDD VDD X3_NET12 X3_NET14  SKY130_FD_SC_HD__FA_1
*--------END___X3_X76->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X77->SKY130_FD_SC_HD__FA_1
X77_X3 RAW_BIT11 RAW_BIT8 RAW_BIT12 VSS VSS VDD VDD X3_NET13 X3_NET15  SKY130_FD_SC_HD__FA_1
*--------END___X3_X77->SKY130_FD_SC_HD__FA_1
*--------BEGIN_X3_X78->SKY130_FD_SC_HD__DFRTP_1
X78_X3 CYCLE31 X3_NET14 RESET VSS VSS VDD VDD BIT8  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X78->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X79->SKY130_FD_SC_HD__DFRTP_1
X79_X3 CYCLE31 X3_NET15 RESET VSS VSS VDD VDD BIT9  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X79->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X80->SKY130_FD_SC_HD__DFRTP_1
X80_X3 CYCLE31 X3_NET16 RESET VSS VSS VDD VDD BIT1  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X80->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X81->SKY130_FD_SC_HD__DFRTP_1
X81_X3 CYCLE31 RAW_BIT13 RESET VSS VSS VDD VDD BIT10  SKY130_FD_SC_HD__DFRTP_1
*--------END___X3_X81->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X3_X82->SKY130_FD_SC_HD__INV_1
X82_X3 CYCLE31 VSS VSS VDD VDD DONE  SKY130_FD_SC_HD__INV_1
*--------END___X3_X82->SKY130_FD_SC_HD__INV_1
*--------END___X3->DEC
*--------BEGIN_X4->RAW_BIT_CALCULATOR
*.PININFO CYCLE[13..1]:I SW_N_SP[9..1]:O VSS:B VDD:B SW_N[8..1]:O SW_P_SP[9..1]:O SW_P[8..1]:O
*+ VCMP:I RESET:I RAW_BIT[13..1]:O
*--------BEGIN_X4_X29->SKY130_FD_SC_HD__XOR2_1
X29_X4 RAW_BIT1 VCMP VSS VSS VDD VDD X4_NET50  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X29->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X31->SKY130_FD_SC_HD__XOR2_1
X31_X4 RAW_BIT1 VCMP VSS VSS VDD VDD X4_NET51  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X31->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X37->SKY130_FD_SC_HD__XOR2_1
X37_X4 RAW_BIT4 VCMP VSS VSS VDD VDD X4_NET52  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X37->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X40->SKY130_FD_SC_HD__XOR2_1
X40_X4 RAW_BIT4 VCMP VSS VSS VDD VDD X4_NET53  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X40->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X45->SKY130_FD_SC_HD__XOR2_1
X45_X4 RAW_BIT4 VCMP VSS VSS VDD VDD X4_NET54  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X45->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X100->SKY130_FD_SC_HD__DFRTP_1
X100_X4 CYCLE18 X4_NET10 X4_NET22 VSS VSS VDD VDD SW_P_SP1  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X100->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X99->SKY130_FD_SC_HD__INV_1
X99_X4 VCMP VSS VSS VDD VDD X4_NET10  SKY130_FD_SC_HD__INV_1
*--------END___X4_X99->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X102->SKY130_FD_SC_HD__DFRTP_1
X102_X4 CYCLE18 VCMP X4_NET22 VSS VSS VDD VDD SW_N_SP1  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X102->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X25->SKY130_FD_SC_HD__DFRTP_1
X25_X4 CYCLE18 VCMP X4_NET24 VSS VSS VDD VDD SW_N_SP2  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X25->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X103->SKY130_FD_SC_HD__INV_1
X103_X4 VCMP VSS VSS VDD VDD X4_NET11  SKY130_FD_SC_HD__INV_1
*--------END___X4_X103->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X104->SKY130_FD_SC_HD__DFRTP_1
X104_X4 CYCLE18 X4_NET11 X4_NET24 VSS VSS VDD VDD SW_P_SP2  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X104->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X21->SKY130_FD_SC_HD__DFSTP_1
X21_X4 X4_NET1 VCMP NET1 VSS VSS VDD VDD SW_N1  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X21->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X22->SKY130_FD_SC_HD__DFSTP_1
X22_X4 X4_NET1 X4_NET12 NET1 VSS VSS VDD VDD SW_P1  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X22->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X105->SKY130_FD_SC_HD__INV_1
X105_X4 VCMP VSS VSS VDD VDD X4_NET12  SKY130_FD_SC_HD__INV_1
*--------END___X4_X105->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X28->SKY130_FD_SC_HD__DFSTP_1
X28_X4 X4_NET3 VCMP NET1 VSS VSS VDD VDD SW_N2  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X28->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X106->SKY130_FD_SC_HD__DFSTP_1
X106_X4 X4_NET3 X4_NET13 NET1 VSS VSS VDD VDD SW_P2  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X106->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X107->SKY130_FD_SC_HD__INV_1
X107_X4 VCMP VSS VSS VDD VDD X4_NET13  SKY130_FD_SC_HD__INV_1
*--------END___X4_X107->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X109->SKY130_FD_SC_HD__INV_1
X109_X4 VCMP VSS VSS VDD VDD X4_NET14  SKY130_FD_SC_HD__INV_1
*--------END___X4_X109->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X111->SKY130_FD_SC_HD__INV_1
X111_X4 VCMP VSS VSS VDD VDD X4_NET15  SKY130_FD_SC_HD__INV_1
*--------END___X4_X111->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X27->SKY130_FD_SC_HD__DFRTP_1
X27_X4 CYCLE21 VCMP X4_NET26 VSS VSS VDD VDD SW_N_SP3  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X27->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X35->SKY130_FD_SC_HD__DFRTP_1
X35_X4 CYCLE21 X4_NET14 X4_NET26 VSS VSS VDD VDD SW_P_SP3  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X35->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X41->SKY130_FD_SC_HD__DFRTP_1
X41_X4 CYCLE21 VCMP X4_NET27 VSS VSS VDD VDD SW_N_SP4  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X41->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X108->SKY130_FD_SC_HD__DFRTP_1
X108_X4 CYCLE21 X4_NET15 X4_NET27 VSS VSS VDD VDD SW_P_SP4  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X108->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X110->SKY130_FD_SC_HD__DFRTP_1
X110_X4 CYCLE21 VCMP X4_NET28 VSS VSS VDD VDD SW_N_SP5  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X110->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X112->SKY130_FD_SC_HD__DFRTP_1
X112_X4 CYCLE21 X4_NET16 X4_NET28 VSS VSS VDD VDD SW_P_SP5  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X112->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X113->SKY130_FD_SC_HD__INV_1
X113_X4 VCMP VSS VSS VDD VDD X4_NET16  SKY130_FD_SC_HD__INV_1
*--------END___X4_X113->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X114->SKY130_FD_SC_HD__DFSTP_1
X114_X4 X4_NET5 X4_NET17 NET1 VSS VSS VDD VDD SW_P3  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X114->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X32->SKY130_FD_SC_HD__DFSTP_1
X32_X4 X4_NET5 VCMP NET1 VSS VSS VDD VDD SW_N3  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X32->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X115->SKY130_FD_SC_HD__INV_1
X115_X4 VCMP VSS VSS VDD VDD X4_NET17  SKY130_FD_SC_HD__INV_1
*--------END___X4_X115->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X38->SKY130_FD_SC_HD__DFSTP_1
X38_X4 X4_NET6 VCMP NET1 VSS VSS VDD VDD SW_N4  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X38->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X116->SKY130_FD_SC_HD__DFSTP_1
X116_X4 X4_NET6 X4_NET18 NET1 VSS VSS VDD VDD SW_P4  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X116->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X117->SKY130_FD_SC_HD__INV_1
X117_X4 VCMP VSS VSS VDD VDD X4_NET18  SKY130_FD_SC_HD__INV_1
*--------END___X4_X117->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X43->SKY130_FD_SC_HD__DFSTP_1
X43_X4 X4_NET7 VCMP NET1 VSS VSS VDD VDD SW_N5  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X43->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X118->SKY130_FD_SC_HD__DFSTP_1
X118_X4 X4_NET7 X4_NET19 NET1 VSS VSS VDD VDD SW_P5  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X118->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X119->SKY130_FD_SC_HD__INV_1
X119_X4 VCMP VSS VSS VDD VDD X4_NET19  SKY130_FD_SC_HD__INV_1
*--------END___X4_X119->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X132->SKY130_FD_SC_HD__DFRTP_1
X132_X4 CYCLE29 X4_NET20 NET1 VSS VSS VDD VDD SW_P_SP9  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X132->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X133->SKY130_FD_SC_HD__INV_1
X133_X4 VCMP VSS VSS VDD VDD X4_NET20  SKY130_FD_SC_HD__INV_1
*--------END___X4_X133->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X61->SKY130_FD_SC_HD__DFRTP_1
X61_X4 CYCLE29 VCMP NET1 VSS VSS VDD VDD SW_N_SP9  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X61->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X24->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X24_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X24 X4_X24_NET1 CYCLE19 VSS VSS VDD VDD X4_NET1  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X24_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X24_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X24 X4_NET50 CYCLE19 VSS VSS VDD VDD X4_NET2  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X24_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X24_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X24 X4_NET50 VSS VSS VDD VDD X4_X24_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X24_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X24->DEMUX2
*--------BEGIN_X4_X30->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X30_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X30 X4_X30_NET1 CYCLE20 VSS VSS VDD VDD X4_NET3  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X30_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X30_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X30 X4_NET51 CYCLE20 VSS VSS VDD VDD X4_NET4  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X30_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X30_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X30 X4_NET51 VSS VSS VDD VDD X4_X30_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X30_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X30->DEMUX2
*--------BEGIN_X4_X34->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X34_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X34 X4_X34_NET1 CYCLE22 VSS VSS VDD VDD X4_NET5  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X34_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X34_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X34 X4_NET52 CYCLE22 VSS VSS VDD VDD X4_NET21  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X34_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X34_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X34 X4_NET52 VSS VSS VDD VDD X4_X34_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X34_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X34->DEMUX2
*--------BEGIN_X4_X39->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X39_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X39 X4_X39_NET1 CYCLE23 VSS VSS VDD VDD X4_NET6  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X39_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X39_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X39 X4_NET53 CYCLE23 VSS VSS VDD VDD X4_NET8  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X39_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X39_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X39 X4_NET53 VSS VSS VDD VDD X4_X39_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X39_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X39->DEMUX2
*--------BEGIN_X4_X44->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X44_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X44 X4_X44_NET1 CYCLE24 VSS VSS VDD VDD X4_NET7  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X44_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X44_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X44 X4_NET54 CYCLE24 VSS VSS VDD VDD X4_NET9  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X44_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X44_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X44 X4_NET54 VSS VSS VDD VDD X4_X44_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X44_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X44->DEMUX2
*--------BEGIN_X4_X1->SKY130_FD_SC_HD__INV_1
X1_X4 X4_NET2 VSS VSS VDD VDD X4_NET23  SKY130_FD_SC_HD__INV_1
*--------END___X4_X1->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X2->SKY130_FD_SC_HD__INV_1
X2_X4 X4_NET4 VSS VSS VDD VDD X4_NET25  SKY130_FD_SC_HD__INV_1
*--------END___X4_X2->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X3->SKY130_FD_SC_HD__DFRTP_4
X3_X4 CYCLE18 VCMP NET1 VSS VSS VDD VDD RAW_BIT1  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X3->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X4->SKY130_FD_SC_HD__DFRTP_4
X4_X4 CYCLE19 VCMP NET1 VSS VSS VDD VDD RAW_BIT2  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X4->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X5->SKY130_FD_SC_HD__DFRTP_4
X5_X4 CYCLE20 VCMP NET1 VSS VSS VDD VDD RAW_BIT3  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X5->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X6->SKY130_FD_SC_HD__DFRTP_4
X6_X4 CYCLE21 VCMP NET1 VSS VSS VDD VDD RAW_BIT4  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X6->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X7->SKY130_FD_SC_HD__DFRTP_4
X7_X4 CYCLE22 VCMP NET1 VSS VSS VDD VDD RAW_BIT5  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X7->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X8->SKY130_FD_SC_HD__DFRTP_4
X8_X4 CYCLE23 VCMP NET1 VSS VSS VDD VDD RAW_BIT6  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X8->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X9->SKY130_FD_SC_HD__DFRTP_4
X9_X4 CYCLE24 VCMP NET1 VSS VSS VDD VDD RAW_BIT7  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X9->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X10->SKY130_FD_SC_HD__DFRTP_4
X10_X4 CYCLE25 VCMP NET1 VSS VSS VDD VDD RAW_BIT8  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X10->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X11->SKY130_FD_SC_HD__DFRTP_4
X11_X4 CYCLE26 VCMP NET1 VSS VSS VDD VDD RAW_BIT9  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X11->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X12->SKY130_FD_SC_HD__DFRTP_4
X12_X4 CYCLE27 VCMP NET1 VSS VSS VDD VDD RAW_BIT10  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X12->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X13->SKY130_FD_SC_HD__DFRTP_4
X13_X4 CYCLE28 VCMP NET1 VSS VSS VDD VDD RAW_BIT11  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X13->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X14->SKY130_FD_SC_HD__DFRTP_4
X14_X4 CYCLE29 VCMP NET1 VSS VSS VDD VDD RAW_BIT12  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X14->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X15->SKY130_FD_SC_HD__DFRTP_4
X15_X4 CYCLE30 VCMP NET1 VSS VSS VDD VDD RAW_BIT13  SKY130_FD_SC_HD__DFRTP_4
*--------END___X4_X15->SKY130_FD_SC_HD__DFRTP_4
*--------BEGIN_X4_X18->SKY130_FD_SC_HD__INV_1
X18_X4 X4_NET21 VSS VSS VDD VDD X4_NET29  SKY130_FD_SC_HD__INV_1
*--------END___X4_X18->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X19->SKY130_FD_SC_HD__INV_1
X19_X4 X4_NET8 VSS VSS VDD VDD X4_NET30  SKY130_FD_SC_HD__INV_1
*--------END___X4_X19->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X20->SKY130_FD_SC_HD__INV_1
X20_X4 X4_NET9 VSS VSS VDD VDD X4_NET31  SKY130_FD_SC_HD__INV_1
*--------END___X4_X20->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X42->SKY130_FD_SC_HD__XOR2_1
X42_X4 RAW_BIT8 VCMP VSS VSS VDD VDD X4_NET55  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X42->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X62->SKY130_FD_SC_HD__XOR2_1
X62_X4 RAW_BIT8 VCMP VSS VSS VDD VDD X4_NET56  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X62->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X64->SKY130_FD_SC_HD__XOR2_1
X64_X4 RAW_BIT8 VCMP VSS VSS VDD VDD X4_NET57  SKY130_FD_SC_HD__XOR2_1
*--------END___X4_X64->SKY130_FD_SC_HD__XOR2_1
*--------BEGIN_X4_X65->SKY130_FD_SC_HD__INV_1
X65_X4 VCMP VSS VSS VDD VDD X4_NET37  SKY130_FD_SC_HD__INV_1
*--------END___X4_X65->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X66->SKY130_FD_SC_HD__INV_1
X66_X4 VCMP VSS VSS VDD VDD X4_NET38  SKY130_FD_SC_HD__INV_1
*--------END___X4_X66->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X67->SKY130_FD_SC_HD__DFRTP_1
X67_X4 CYCLE25 VCMP X4_NET44 VSS VSS VDD VDD SW_N_SP6  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X67->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X68->SKY130_FD_SC_HD__DFRTP_1
X68_X4 CYCLE25 X4_NET37 X4_NET44 VSS VSS VDD VDD SW_P_SP6  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X68->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X69->SKY130_FD_SC_HD__DFRTP_1
X69_X4 CYCLE25 VCMP X4_NET45 VSS VSS VDD VDD SW_N_SP7  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X69->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X70->SKY130_FD_SC_HD__DFRTP_1
X70_X4 CYCLE25 X4_NET38 X4_NET45 VSS VSS VDD VDD SW_P_SP7  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X70->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X71->SKY130_FD_SC_HD__DFRTP_1
X71_X4 CYCLE25 VCMP X4_NET46 VSS VSS VDD VDD SW_N_SP8  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X71->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X72->SKY130_FD_SC_HD__DFRTP_1
X72_X4 CYCLE25 X4_NET39 X4_NET46 VSS VSS VDD VDD SW_P_SP8  SKY130_FD_SC_HD__DFRTP_1
*--------END___X4_X72->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X4_X73->SKY130_FD_SC_HD__INV_1
X73_X4 VCMP VSS VSS VDD VDD X4_NET39  SKY130_FD_SC_HD__INV_1
*--------END___X4_X73->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X74->SKY130_FD_SC_HD__DFSTP_1
X74_X4 X4_NET32 X4_NET40 NET1 VSS VSS VDD VDD SW_P6  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X74->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X75->SKY130_FD_SC_HD__DFSTP_1
X75_X4 X4_NET32 VCMP NET1 VSS VSS VDD VDD SW_N6  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X75->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X76->SKY130_FD_SC_HD__INV_1
X76_X4 VCMP VSS VSS VDD VDD X4_NET40  SKY130_FD_SC_HD__INV_1
*--------END___X4_X76->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X77->SKY130_FD_SC_HD__DFSTP_1
X77_X4 X4_NET33 VCMP NET1 VSS VSS VDD VDD SW_N7  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X77->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X78->SKY130_FD_SC_HD__DFSTP_1
X78_X4 X4_NET33 X4_NET41 NET1 VSS VSS VDD VDD SW_P7  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X78->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X79->SKY130_FD_SC_HD__INV_1
X79_X4 VCMP VSS VSS VDD VDD X4_NET41  SKY130_FD_SC_HD__INV_1
*--------END___X4_X79->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X80->SKY130_FD_SC_HD__DFSTP_1
X80_X4 X4_NET34 VCMP NET1 VSS VSS VDD VDD SW_N8  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X80->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X81->SKY130_FD_SC_HD__DFSTP_1
X81_X4 X4_NET34 X4_NET42 NET1 VSS VSS VDD VDD SW_P8  SKY130_FD_SC_HD__DFSTP_1
*--------END___X4_X81->SKY130_FD_SC_HD__DFSTP_1
*--------BEGIN_X4_X82->SKY130_FD_SC_HD__INV_1
X82_X4 VCMP VSS VSS VDD VDD X4_NET42  SKY130_FD_SC_HD__INV_1
*--------END___X4_X82->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X83->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X83_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X83 X4_X83_NET1 CYCLE26 VSS VSS VDD VDD X4_NET32  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X83_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X83_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X83 X4_NET55 CYCLE26 VSS VSS VDD VDD X4_NET43  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X83_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X83_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X83 X4_NET55 VSS VSS VDD VDD X4_X83_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X83_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X83->DEMUX2
*--------BEGIN_X4_X84->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X84_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X84 X4_X84_NET1 CYCLE27 VSS VSS VDD VDD X4_NET33  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X84_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X84_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X84 X4_NET56 CYCLE27 VSS VSS VDD VDD X4_NET35  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X84_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X84_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X84 X4_NET56 VSS VSS VDD VDD X4_X84_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X84_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X84->DEMUX2
*--------BEGIN_X4_X85->DEMUX2
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
*--------BEGIN_X4_X85_X1->SKY130_FD_SC_HD__AND2_0
X1_X4_X85 X4_X85_NET1 CYCLE28 VSS VSS VDD VDD X4_NET34  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X85_X1->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X85_X2->SKY130_FD_SC_HD__AND2_0
X2_X4_X85 X4_NET57 CYCLE28 VSS VSS VDD VDD X4_NET36  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X85_X2->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X85_X3->SKY130_FD_SC_HD__INV_1
X3_X4_X85 X4_NET57 VSS VSS VDD VDD X4_X85_NET1  SKY130_FD_SC_HD__INV_1
*--------END___X4_X85_X3->SKY130_FD_SC_HD__INV_1
*--------END___X4_X85->DEMUX2
*--------BEGIN_X4_X88->SKY130_FD_SC_HD__INV_1
X88_X4 X4_NET43 VSS VSS VDD VDD X4_NET47  SKY130_FD_SC_HD__INV_1
*--------END___X4_X88->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X89->SKY130_FD_SC_HD__INV_1
X89_X4 X4_NET35 VSS VSS VDD VDD X4_NET48  SKY130_FD_SC_HD__INV_1
*--------END___X4_X89->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X90->SKY130_FD_SC_HD__INV_1
X90_X4 X4_NET36 VSS VSS VDD VDD X4_NET49  SKY130_FD_SC_HD__INV_1
*--------END___X4_X90->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X4_X46->SKY130_FD_SC_HD__AND2_0
X46_X4 X4_NET23 NET1 VSS VSS VDD VDD X4_NET22  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X46->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X23->SKY130_FD_SC_HD__AND2_0
X23_X4 X4_NET25 NET1 VSS VSS VDD VDD X4_NET24  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X23->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X26->SKY130_FD_SC_HD__AND2_0
X26_X4 X4_NET29 NET1 VSS VSS VDD VDD X4_NET26  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X26->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X16->SKY130_FD_SC_HD__AND2_0
X16_X4 X4_NET30 NET1 VSS VSS VDD VDD X4_NET27  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X16->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X17->SKY130_FD_SC_HD__AND2_0
X17_X4 X4_NET31 NET1 VSS VSS VDD VDD X4_NET28  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X17->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X33->SKY130_FD_SC_HD__AND2_0
X33_X4 X4_NET47 NET1 VSS VSS VDD VDD X4_NET44  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X33->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X36->SKY130_FD_SC_HD__AND2_0
X36_X4 X4_NET48 NET1 VSS VSS VDD VDD X4_NET45  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X36->SKY130_FD_SC_HD__AND2_0
*--------BEGIN_X4_X47->SKY130_FD_SC_HD__AND2_0
X47_X4 X4_NET49 NET1 VSS VSS VDD VDD X4_NET46  SKY130_FD_SC_HD__AND2_0
*--------END___X4_X47->SKY130_FD_SC_HD__AND2_0
*--------END___X4->RAW_BIT_CALCULATOR
*--------BEGIN_X1->SHIFTED_CLOCK_GENERATOR
*.PININFO CYCLE[31..0]:O VSS:B VDD:B CLK:I RESET:I
*--------BEGIN_X1_X32->SKY130_FD_SC_HD__DFRTP_1
X32_X1 CLK CYCLE0 X1_RESET_B VSS VSS VDD VDD CYCLE1  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X32->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X1->SKY130_FD_SC_HD__DFRTP_1
X1_X1 CLK CYCLE1 X1_RESET_B VSS VSS VDD VDD CYCLE2  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X1->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X2->SKY130_FD_SC_HD__DFRTP_1
X2_X1 CLK CYCLE2 X1_RESET_B VSS VSS VDD VDD CYCLE3  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X2->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X3->SKY130_FD_SC_HD__DFRTP_1
X3_X1 CLK CYCLE3 X1_RESET_B VSS VSS VDD VDD CYCLE4  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X3->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X4->SKY130_FD_SC_HD__DFRTP_1
X4_X1 CLK CYCLE4 X1_RESET_B VSS VSS VDD VDD CYCLE5  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X4->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X5->SKY130_FD_SC_HD__DFRTP_1
X5_X1 CLK CYCLE5 X1_RESET_B VSS VSS VDD VDD CYCLE6  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X5->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X6->SKY130_FD_SC_HD__DFRTP_1
X6_X1 CLK CYCLE6 X1_RESET_B VSS VSS VDD VDD CYCLE7  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X6->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X7->SKY130_FD_SC_HD__DFRTP_1
X7_X1 CLK CYCLE7 X1_RESET_B VSS VSS VDD VDD CYCLE8  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X7->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X8->SKY130_FD_SC_HD__DFRTP_1
X8_X1 CLK CYCLE8 X1_RESET_B VSS VSS VDD VDD CYCLE9  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X8->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X9->SKY130_FD_SC_HD__DFRTP_1
X9_X1 CLK CYCLE9 X1_RESET_B VSS VSS VDD VDD CYCLE10  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X9->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X10->SKY130_FD_SC_HD__DFRTP_1
X10_X1 CLK CYCLE10 X1_RESET_B VSS VSS VDD VDD CYCLE11  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X10->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X11->SKY130_FD_SC_HD__DFRTP_1
X11_X1 CLK CYCLE11 X1_RESET_B VSS VSS VDD VDD CYCLE12  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X11->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X12->SKY130_FD_SC_HD__DFRTP_1
X12_X1 CLK CYCLE12 X1_RESET_B VSS VSS VDD VDD CYCLE13  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X12->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X13->SKY130_FD_SC_HD__DFRTP_1
X13_X1 CLK CYCLE13 X1_RESET_B VSS VSS VDD VDD CYCLE14  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X13->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X14->SKY130_FD_SC_HD__DFRTP_1
X14_X1 CLK CYCLE14 X1_RESET_B VSS VSS VDD VDD CYCLE15  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X14->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X15->SKY130_FD_SC_HD__DFRTP_1
X15_X1 CLK CYCLE15 X1_RESET_B VSS VSS VDD VDD CYCLE16  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X15->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X16->SKY130_FD_SC_HD__DFRTP_1
X16_X1 CLK CYCLE16 X1_RESET_B VSS VSS VDD VDD CYCLE17  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X16->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X17->SKY130_FD_SC_HD__DFRTP_1
X17_X1 CLK CYCLE17 X1_RESET_B VSS VSS VDD VDD CYCLE18  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X17->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X18->SKY130_FD_SC_HD__DFRTP_1
X18_X1 CLK CYCLE18 X1_RESET_B VSS VSS VDD VDD CYCLE19  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X18->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X19->SKY130_FD_SC_HD__DFRTP_1
X19_X1 CLK CYCLE19 X1_RESET_B VSS VSS VDD VDD CYCLE20  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X19->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X20->SKY130_FD_SC_HD__DFRTP_1
X20_X1 CLK CYCLE20 X1_RESET_B VSS VSS VDD VDD CYCLE21  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X20->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X21->SKY130_FD_SC_HD__DFRTP_1
X21_X1 CLK CYCLE21 X1_RESET_B VSS VSS VDD VDD CYCLE22  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X21->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X22->SKY130_FD_SC_HD__DFRTP_1
X22_X1 CLK CYCLE22 X1_RESET_B VSS VSS VDD VDD CYCLE23  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X22->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X23->SKY130_FD_SC_HD__DFRTP_1
X23_X1 CLK CYCLE23 X1_RESET_B VSS VSS VDD VDD CYCLE24  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X23->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X24->SKY130_FD_SC_HD__DFRTP_1
X24_X1 CLK CYCLE24 X1_RESET_B VSS VSS VDD VDD CYCLE25  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X24->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X25->SKY130_FD_SC_HD__DFRTP_1
X25_X1 CLK CYCLE25 X1_RESET_B VSS VSS VDD VDD CYCLE26  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X25->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X26->SKY130_FD_SC_HD__DFRTP_1
X26_X1 CLK CYCLE26 X1_RESET_B VSS VSS VDD VDD CYCLE27  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X26->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X27->SKY130_FD_SC_HD__DFRTP_1
X27_X1 CLK CYCLE27 X1_RESET_B VSS VSS VDD VDD CYCLE28  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X27->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X28->SKY130_FD_SC_HD__DFRTP_1
X28_X1 CLK CYCLE28 X1_RESET_B VSS VSS VDD VDD CYCLE29  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X28->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X29->SKY130_FD_SC_HD__DFRTP_1
X29_X1 CLK CYCLE29 X1_RESET_B VSS VSS VDD VDD CYCLE30  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X29->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X30->SKY130_FD_SC_HD__DFRTP_1
X30_X1 CLK CYCLE30 X1_RESET_B VSS VSS VDD VDD CYCLE31  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X30->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X31->SKY130_FD_SC_HD__DFRTP_1
X31_X1 CLK VDD X1_RESET_B VSS VSS VDD VDD CYCLE0  SKY130_FD_SC_HD__DFRTP_1
*--------END___X1_X31->SKY130_FD_SC_HD__DFRTP_1
*--------BEGIN_X1_X37->SKY130_FD_SC_HD__BUF_16
X37_X1 X1_NET1 VSS VSS VDD VDD X1_RESET_B  SKY130_FD_SC_HD__BUF_16
*--------END___X1_X37->SKY130_FD_SC_HD__BUF_16
*--------BEGIN_X1_X35->SKY130_FD_SC_HD__AND2_4
X35_X1 X1_RESET_CYCLE RESET VSS VSS VDD VDD X1_NET1  SKY130_FD_SC_HD__AND2_4
*--------END___X1_X35->SKY130_FD_SC_HD__AND2_4
*--------BEGIN_X1_X33->SKY130_FD_SC_HD__DFRTN_1
X33_X1 CLK CYCLE31 X1_RESET_B VSS VSS VDD VDD X1_HALF_CYCLE  SKY130_FD_SC_HD__DFRTN_1
*--------END___X1_X33->SKY130_FD_SC_HD__DFRTN_1
*--------BEGIN_X1_X38->SKY130_FD_SC_HD__NAND2_1
X38_X1 X1_HALF_CYCLE CYCLE31 VSS VSS VDD VDD X1_RESET_CYCLE  SKY130_FD_SC_HD__NAND2_1
*--------END___X1_X38->SKY130_FD_SC_HD__NAND2_1
*--------END___X1->SHIFTED_CLOCK_GENERATOR
*--------BEGIN_X8->SKY130_FD_SC_HD__OR4_2
X8 NET2 NET3 NET5 NET4 VSS VSS VDD VDD NET6  SKY130_FD_SC_HD__OR4_2
*--------END___X8->SKY130_FD_SC_HD__OR4_2
*--------BEGIN_X9->SKY130_FD_SC_HD__DFRTN_1
X9 CLK NET6 RESET VSS VSS VDD VDD SW_SAMPLE  SKY130_FD_SC_HD__DFRTN_1
*--------END___X9->SKY130_FD_SC_HD__DFRTN_1
*--------BEGIN_X10->SKY130_FD_SC_HD__OR3_2
X10 CYCLE13 CYCLE14 CYCLE15 VSS VSS VDD VDD NET4  SKY130_FD_SC_HD__OR3_2
*--------END___X10->SKY130_FD_SC_HD__OR3_2
*--------BEGIN_X6->SKY130_FD_SC_HD__INV_16
X6 CYCLE0 VSS VSS VDD VDD NET1  SKY130_FD_SC_HD__INV_16
*--------END___X6->SKY130_FD_SC_HD__INV_16
.end
