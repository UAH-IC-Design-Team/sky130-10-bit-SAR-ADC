magic
tech sky130A
magscale 1 2
timestamp 1666555793
<< checkpaint >>
rect 7569 7901 10511 31638
rect -153 7323 10511 7901
rect 17872 7323 20814 31060
rect -153 2514 20814 7323
rect -944 1807 20814 2514
rect -944 1354 21183 1807
rect -944 -766 21552 1354
rect -575 -819 21552 -766
rect 6093 -872 21552 -819
rect 6462 -925 21552 -872
rect 6831 -978 21552 -925
rect 7200 -1031 21552 -978
rect 7569 -1084 21552 -1031
rect 7938 -1137 21552 -1084
rect 8307 -1190 21552 -1137
rect 9359 -1344 21552 -1190
rect 9728 -1397 21552 -1344
rect 16396 -1450 21552 -1397
rect 16765 -1503 21552 -1450
rect 17134 -1556 21552 -1503
rect 17503 -1609 21552 -1556
rect 17872 -1662 21552 -1609
rect 18241 -1715 21552 -1662
rect 18610 -1768 21552 -1715
<< error_s >>
rect 9011 5148 9069 5154
rect 9011 5114 9023 5148
rect 9011 5108 9069 5114
rect 9011 5040 9069 5046
rect 9011 5006 9023 5040
rect 9011 5000 9069 5006
rect 9011 4748 9069 4754
rect 9011 4714 9023 4748
rect 9011 4708 9069 4714
rect 9011 4640 9069 4646
rect 9011 4606 9023 4640
rect 9011 4600 9069 4606
rect 9011 4348 9069 4354
rect 9011 4314 9023 4348
rect 9011 4308 9069 4314
rect 9011 4240 9069 4246
rect 9011 4206 9023 4240
rect 9011 4200 9069 4206
rect 9011 3948 9069 3954
rect 9011 3914 9023 3948
rect 9011 3908 9069 3914
rect 9011 3840 9069 3846
rect 129 3811 187 3817
rect 129 3777 141 3811
rect 9011 3806 9023 3840
rect 9011 3800 9069 3806
rect 129 3771 187 3777
rect 9011 3548 9069 3554
rect 129 3519 187 3525
rect 129 3485 141 3519
rect 9011 3514 9023 3548
rect 9011 3508 9069 3514
rect 129 3479 187 3485
rect 9011 3440 9069 3446
rect 129 3411 187 3417
rect 129 3377 141 3411
rect 9011 3406 9023 3440
rect 9011 3400 9069 3406
rect 129 3371 187 3377
rect 10432 3233 10490 3239
rect 10432 3199 10444 3233
rect 10432 3193 10490 3199
rect 9011 3148 9069 3154
rect 129 3119 187 3125
rect 129 3085 141 3119
rect 9011 3114 9023 3148
rect 9011 3108 9069 3114
rect 129 3079 187 3085
rect 9011 3040 9069 3046
rect 129 3011 187 3017
rect 129 2977 141 3011
rect 9011 3006 9023 3040
rect 9011 3000 9069 3006
rect 129 2971 187 2977
rect 10432 2941 10490 2947
rect 10432 2907 10444 2941
rect 10432 2901 10490 2907
rect 10432 2833 10490 2839
rect 10432 2799 10444 2833
rect 10432 2793 10490 2799
rect 9011 2748 9069 2754
rect 129 2719 187 2725
rect 129 2685 141 2719
rect 9011 2714 9023 2748
rect 9011 2708 9069 2714
rect 129 2679 187 2685
rect 9011 2640 9069 2646
rect 129 2611 187 2617
rect 129 2577 141 2611
rect 9011 2606 9023 2640
rect 9011 2600 9069 2606
rect 129 2571 187 2577
rect 10432 2541 10490 2547
rect 10432 2507 10444 2541
rect 10432 2501 10490 2507
rect 10432 2433 10490 2439
rect 10432 2399 10444 2433
rect 10432 2393 10490 2399
rect 9011 2348 9069 2354
rect 129 2319 187 2325
rect 129 2285 141 2319
rect 9011 2314 9023 2348
rect 9011 2308 9069 2314
rect 129 2279 187 2285
rect 9011 2240 9069 2246
rect 129 2211 187 2217
rect 129 2177 141 2211
rect 9011 2206 9023 2240
rect 9011 2200 9069 2206
rect 129 2171 187 2177
rect 10432 2141 10490 2147
rect 10432 2107 10444 2141
rect 10432 2101 10490 2107
rect 10432 2033 10490 2039
rect 10432 1999 10444 2033
rect 10432 1993 10490 1999
rect 9011 1948 9069 1954
rect 129 1919 187 1925
rect 129 1885 141 1919
rect 9011 1914 9023 1948
rect 9011 1908 9069 1914
rect 129 1879 187 1885
rect 9011 1840 9069 1846
rect 129 1811 187 1817
rect 129 1777 141 1811
rect 9011 1806 9023 1840
rect 9011 1800 9069 1806
rect 129 1771 187 1777
rect 10432 1741 10490 1747
rect 10432 1707 10444 1741
rect 10432 1701 10490 1707
rect 7535 1688 7593 1694
rect 7535 1654 7547 1688
rect 7535 1648 7593 1654
rect 10432 1633 10490 1639
rect 10432 1599 10444 1633
rect 10432 1593 10490 1599
rect 9011 1548 9069 1554
rect 129 1519 187 1525
rect 129 1485 141 1519
rect 9011 1514 9023 1548
rect 9011 1508 9069 1514
rect 129 1479 187 1485
rect 9011 1440 9069 1446
rect 129 1411 187 1417
rect 129 1377 141 1411
rect 9011 1406 9023 1440
rect 9011 1400 9069 1406
rect 129 1371 187 1377
rect 10432 1341 10490 1347
rect 10432 1307 10444 1341
rect 10432 1301 10490 1307
rect 299 1254 333 1272
rect 299 1218 369 1254
rect 10432 1233 10490 1239
rect 316 1184 387 1218
rect 10432 1199 10444 1233
rect 10432 1193 10490 1199
rect 129 1119 187 1125
rect 129 1085 141 1119
rect 129 1079 187 1085
rect 129 1011 187 1017
rect 129 977 141 1011
rect 129 971 187 977
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1184
rect 9011 1148 9069 1154
rect 498 1116 556 1122
rect 498 1082 510 1116
rect 9011 1114 9023 1148
rect 498 1076 556 1082
rect 668 1043 702 1061
rect 7705 1059 7739 1113
rect 9011 1108 9069 1114
rect 9181 1089 9215 1143
rect 668 1007 738 1043
rect 685 973 756 1007
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 685 530 755 973
rect 867 905 925 911
rect 867 871 879 905
rect 867 865 925 871
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 7535 560 7593 566
rect 685 494 738 530
rect 7535 526 7547 560
rect 7535 520 7593 526
rect 7724 424 7739 1059
rect 7758 1025 7793 1059
rect 9011 1040 9069 1046
rect 7758 424 7792 1025
rect 9011 1006 9023 1040
rect 9011 1000 9069 1006
rect 7904 957 7962 963
rect 7904 923 7916 957
rect 7904 917 7962 923
rect 8074 884 8108 902
rect 8074 848 8144 884
rect 8091 814 8162 848
rect 8442 814 8477 848
rect 7904 507 7962 513
rect 7904 473 7916 507
rect 7904 467 7962 473
rect 7758 390 7773 424
rect 8091 371 8161 814
rect 8443 795 8477 814
rect 8273 746 8331 752
rect 8273 712 8285 746
rect 8273 706 8331 712
rect 8273 454 8331 460
rect 8273 420 8285 454
rect 8273 414 8331 420
rect 8091 335 8144 371
rect 8462 318 8477 795
rect 8496 761 8531 795
rect 8496 318 8530 761
rect 8642 693 8700 699
rect 8642 659 8654 693
rect 8642 653 8700 659
rect 8642 401 8700 407
rect 8642 367 8654 401
rect 8642 361 8700 367
rect 8496 284 8511 318
rect 8831 265 8846 795
rect 8865 265 8899 849
rect 9011 748 9069 754
rect 9011 714 9023 748
rect 9011 708 9069 714
rect 9011 640 9069 646
rect 9011 606 9023 640
rect 9011 600 9069 606
rect 9011 348 9069 354
rect 9011 314 9023 348
rect 9011 308 9069 314
rect 8865 231 8880 265
rect 9200 212 9215 1089
rect 9234 1055 9269 1089
rect 9234 212 9268 1055
rect 9380 987 9438 993
rect 9380 953 9392 987
rect 9380 947 9438 953
rect 10432 941 10490 947
rect 10432 907 10444 941
rect 10432 901 10490 907
rect 10432 833 10490 839
rect 10432 799 10444 833
rect 10432 793 10490 799
rect 9380 695 9438 701
rect 9380 661 9392 695
rect 9380 655 9438 661
rect 9550 636 9584 690
rect 10602 676 10636 694
rect 10286 652 10299 665
rect 9380 587 9438 593
rect 9380 553 9392 587
rect 9380 547 9438 553
rect 9380 295 9438 301
rect 9380 261 9392 295
rect 9380 255 9438 261
rect 9234 178 9249 212
rect 9569 159 9584 636
rect 9603 602 9638 636
rect 9603 159 9637 602
rect 9749 534 9807 540
rect 9749 500 9761 534
rect 9749 494 9807 500
rect 9951 331 9989 652
rect 10250 331 10303 652
rect 10602 640 10672 676
rect 10619 606 10690 640
rect 10432 541 10490 547
rect 10432 507 10444 541
rect 10432 501 10490 507
rect 10432 433 10490 439
rect 10432 399 10444 433
rect 10432 393 10490 399
rect 9749 242 9807 248
rect 9749 208 9761 242
rect 9749 202 9807 208
rect 9603 125 9618 159
rect 10286 121 10292 255
rect 10432 141 10490 147
rect 10252 53 10265 87
rect 10286 19 10299 121
rect 10432 107 10444 141
rect 10432 101 10490 107
rect 10619 5 10689 606
rect 10801 538 10859 544
rect 10801 504 10813 538
rect 10801 498 10859 504
rect 10971 465 11005 483
rect 10971 429 11041 465
rect 10988 395 11059 429
rect 10801 88 10859 94
rect 10801 54 10813 88
rect 10801 48 10859 54
rect 10619 -31 10672 5
rect 10988 -48 11058 395
rect 11170 327 11228 333
rect 11170 293 11182 327
rect 11170 287 11228 293
rect 11170 35 11228 41
rect 11170 1 11182 35
rect 11170 -5 11228 1
rect 10988 -84 11041 -48
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 0
transform 1 0 4257 0 1 3541
box -3150 -3100 3149 3100
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 0
transform 1 0 14560 0 1 2963
box -3150 -3100 3149 3100
use sky130_fd_pr__nfet_01v8_CCZD88  XM1
timestamp 0
transform 1 0 158 0 1 2248
box -211 -1701 211 1701
use sky130_fd_pr__pfet_01v8_NF5F9G  XM2
timestamp 0
transform 1 0 527 0 1 874
box -211 -380 211 380
use sky130_fd_pr__nfet_01v8_77T378  XM3
timestamp 0
transform 1 0 896 0 1 742
box -211 -301 211 301
use sky130_fd_pr__pfet_01v8_UGSVTG  XM4
timestamp 0
transform 1 0 7564 0 1 1107
box -211 -719 211 719
use sky130_fd_pr__pfet_01v8_NF5F9G  XM5
timestamp 0
transform 1 0 7933 0 1 715
box -211 -380 211 380
use sky130_fd_pr__nfet_01v8_77T378  XM6
timestamp 0
transform 1 0 8302 0 1 583
box -211 -301 211 301
use sky130_fd_pr__nfet_01v8_77T378  XM7
timestamp 0
transform 1 0 8671 0 1 530
box -211 -301 211 301
use sky130_fd_pr__nfet_01v8_FBZ6SX  XM8
timestamp 0
transform 1 0 9040 0 1 15277
box -211 -15101 211 15101
use sky130_fd_pr__nfet_01v8_6V4E88  XM9
timestamp 0
transform 1 0 9409 0 1 624
box -211 -501 211 501
use sky130_fd_pr__nfet_01v8_77T378  XM10
timestamp 0
transform 1 0 9778 0 1 371
box -211 -301 211 301
use sky130_fd_pr__nfet_01v8_CCZD88  XM11
timestamp 0
transform 1 0 10461 0 1 1670
box -211 -1701 211 1701
use sky130_fd_pr__pfet_01v8_NF5F9G  XM12
timestamp 0
transform 1 0 10830 0 1 296
box -211 -380 211 380
use sky130_fd_pr__nfet_01v8_77T378  XM13
timestamp 0
transform 1 0 11199 0 1 164
box -211 -301 211 301
use sky130_fd_pr__pfet_01v8_UGSVTG  XM14
timestamp 0
transform 1 0 17867 0 1 529
box -211 -719 211 719
use sky130_fd_pr__pfet_01v8_NF5F9G  XM15
timestamp 0
transform 1 0 18236 0 1 137
box -211 -380 211 380
use sky130_fd_pr__nfet_01v8_77T378  XM16
timestamp 0
transform 1 0 18605 0 1 5
box -211 -301 211 301
use sky130_fd_pr__nfet_01v8_77T378  XM17
timestamp 0
transform 1 0 18974 0 1 -48
box -211 -301 211 301
use sky130_fd_pr__nfet_01v8_FBZ6SX  XM18
timestamp 0
transform 1 0 19343 0 1 14699
box -211 -15101 211 15101
use sky130_fd_pr__nfet_01v8_6V4E88  XM19
timestamp 0
transform 1 0 19712 0 1 46
box -211 -501 211 501
use sky130_fd_pr__nfet_01v8_77T378  XM20
timestamp 0
transform 1 0 20081 0 1 -207
box -211 -301 211 301
use sky130_fd_sc_hd__clkinv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9989 0 1 70
box -38 -48 314 592
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin_p
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout_p
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Vout_n
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Vin_n
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Clk
port 6 nsew
<< end >>
