* NGSPICE file created from demux2.ext - technology: sky130A


* Top level circuit demux2

.end

