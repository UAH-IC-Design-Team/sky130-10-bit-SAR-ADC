magic
tech sky130A
magscale 1 2
timestamp 1665675118
<< error_p >>
rect -70 -2205 -10 2205
rect 10 -2205 70 2205
<< metal3 >>
rect -709 2177 -10 2205
rect -709 -2177 -94 2177
rect -30 -2177 -10 2177
rect -709 -2205 -10 -2177
rect 10 2177 709 2205
rect 10 -2177 625 2177
rect 689 -2177 709 2177
rect 10 -2205 709 -2177
<< via3 >>
rect -94 -2177 -30 2177
rect 625 -2177 689 2177
<< mimcap >>
rect -609 2065 -209 2105
rect -609 -2065 -569 2065
rect -249 -2065 -209 2065
rect -609 -2105 -209 -2065
rect 110 2065 510 2105
rect 110 -2065 150 2065
rect 470 -2065 510 2065
rect 110 -2105 510 -2065
<< mimcapcontact >>
rect -569 -2065 -249 2065
rect 150 -2065 470 2065
<< metal4 >>
rect -110 2177 -14 2193
rect -570 2065 -248 2066
rect -570 -2065 -569 2065
rect -249 -2065 -248 2065
rect -570 -2066 -248 -2065
rect -110 -2177 -94 2177
rect -30 -2177 -14 2177
rect 609 2177 705 2193
rect 149 2065 471 2066
rect 149 -2065 150 2065
rect 470 -2065 471 2065
rect 149 -2066 471 -2065
rect -110 -2193 -14 -2177
rect 609 -2177 625 2177
rect 689 -2177 705 2177
rect 609 -2193 705 -2177
<< properties >>
string FIXED_BBOX 10 -2205 610 2205
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
