magic
tech sky130A
magscale 1 2
timestamp 1666489318
<< error_p >>
rect -407 62 -361 74
rect -215 62 -169 74
rect -23 62 23 74
rect 169 62 215 74
rect 361 62 407 74
rect -407 28 -401 62
rect -215 28 -209 62
rect -23 28 -17 62
rect 169 28 175 62
rect 361 28 367 62
rect -407 16 -361 28
rect -215 16 -169 28
rect -23 16 23 28
rect 169 16 215 28
rect 361 16 407 28
rect -311 -28 -265 -16
rect -119 -28 -73 -16
rect 73 -28 119 -16
rect 265 -28 311 -16
rect -311 -62 -305 -28
rect -119 -62 -113 -28
rect 73 -62 79 -28
rect 265 -62 271 -28
rect -311 -74 -265 -62
rect -119 -74 -73 -62
rect 73 -74 119 -62
rect 265 -74 311 -62
<< nmos >>
rect -351 -91 -321 91
rect -255 -91 -225 91
rect -159 -91 -129 91
rect -63 -91 -33 91
rect 33 -91 63 91
rect 129 -91 159 91
rect 225 -91 255 91
rect 321 -91 351 91
<< ndiff >>
rect -413 79 -351 91
rect -413 -79 -401 79
rect -367 -79 -351 79
rect -413 -91 -351 -79
rect -321 79 -255 91
rect -321 -79 -305 79
rect -271 -79 -255 79
rect -321 -91 -255 -79
rect -225 79 -159 91
rect -225 -79 -209 79
rect -175 -79 -159 79
rect -225 -91 -159 -79
rect -129 79 -63 91
rect -129 -79 -113 79
rect -79 -79 -63 79
rect -129 -91 -63 -79
rect -33 79 33 91
rect -33 -79 -17 79
rect 17 -79 33 79
rect -33 -91 33 -79
rect 63 79 129 91
rect 63 -79 79 79
rect 113 -79 129 79
rect 63 -91 129 -79
rect 159 79 225 91
rect 159 -79 175 79
rect 209 -79 225 79
rect 159 -91 225 -79
rect 255 79 321 91
rect 255 -79 271 79
rect 305 -79 321 79
rect 255 -91 321 -79
rect 351 79 413 91
rect 351 -79 367 79
rect 401 -79 413 79
rect 351 -91 413 -79
<< ndiffc >>
rect -401 -79 -367 79
rect -305 -79 -271 79
rect -209 -79 -175 79
rect -113 -79 -79 79
rect -17 -79 17 79
rect 79 -79 113 79
rect 175 -79 209 79
rect 271 -79 305 79
rect 367 -79 401 79
<< poly >>
rect -351 91 -321 121
rect -255 91 -225 121
rect -159 91 -129 121
rect -63 91 -33 121
rect 33 91 63 121
rect 129 91 159 121
rect 225 91 255 121
rect 321 91 351 121
rect -351 -113 -321 -91
rect -255 -113 -225 -91
rect -159 -113 -129 -91
rect -63 -113 -33 -91
rect 33 -113 63 -91
rect 129 -113 159 -91
rect 225 -113 255 -91
rect 321 -113 351 -91
rect -377 -129 383 -113
rect -377 -163 -353 -129
rect -319 -163 -257 -129
rect -223 -163 -161 -129
rect -127 -163 -67 -129
rect -33 -163 31 -129
rect 65 -163 123 -129
rect 157 -163 223 -129
rect 257 -163 323 -129
rect 357 -163 383 -129
rect -377 -179 383 -163
<< polycont >>
rect -353 -163 -319 -129
rect -257 -163 -223 -129
rect -161 -163 -127 -129
rect -67 -163 -33 -129
rect 31 -163 65 -129
rect 123 -163 157 -129
rect 223 -163 257 -129
rect 323 -163 357 -129
<< locali >>
rect -401 79 -367 95
rect -401 -95 -367 -79
rect -305 79 -271 95
rect -305 -95 -271 -79
rect -209 79 -175 95
rect -209 -95 -175 -79
rect -113 79 -79 95
rect -113 -95 -79 -79
rect -17 79 17 95
rect -17 -95 17 -79
rect 79 79 113 95
rect 79 -95 113 -79
rect 175 79 209 95
rect 175 -95 209 -79
rect 271 79 305 95
rect 271 -95 305 -79
rect 367 79 401 95
rect 367 -95 401 -79
rect -377 -163 -353 -129
rect -319 -163 -257 -129
rect -223 -163 -161 -129
rect -127 -163 -67 -129
rect -33 -163 31 -129
rect 65 -163 123 -129
rect 157 -163 223 -129
rect 257 -163 323 -129
rect 357 -163 383 -129
<< viali >>
rect -401 28 -367 62
rect -305 -62 -271 -28
rect -209 28 -175 62
rect -113 -62 -79 -28
rect -17 28 17 62
rect 79 -62 113 -28
rect 175 28 209 62
rect 271 -62 305 -28
rect 367 28 401 62
rect -353 -163 -319 -129
rect -257 -163 -223 -129
rect -161 -163 -127 -129
rect -67 -163 -33 -129
rect 31 -163 65 -129
rect 123 -163 157 -129
rect 223 -163 257 -129
rect 323 -163 357 -129
<< metal1 >>
rect -407 62 -361 74
rect -407 28 -401 62
rect -367 28 -361 62
rect -407 16 -361 28
rect -215 62 -169 74
rect -215 28 -209 62
rect -175 28 -169 62
rect -215 16 -169 28
rect -23 62 23 74
rect -23 28 -17 62
rect 17 28 23 62
rect -23 16 23 28
rect 169 62 215 74
rect 169 28 175 62
rect 209 28 215 62
rect 169 16 215 28
rect 361 62 407 74
rect 361 28 367 62
rect 401 28 407 62
rect 361 16 407 28
rect -311 -28 -265 -16
rect -311 -62 -305 -28
rect -271 -62 -265 -28
rect -311 -74 -265 -62
rect -119 -28 -73 -16
rect -119 -62 -113 -28
rect -79 -62 -73 -28
rect -119 -74 -73 -62
rect 73 -28 119 -16
rect 73 -62 79 -28
rect 113 -62 119 -28
rect 73 -74 119 -62
rect 265 -28 311 -16
rect 265 -62 271 -28
rect 305 -62 311 -28
rect 265 -74 311 -62
rect -377 -129 383 -123
rect -377 -163 -353 -129
rect -319 -163 -257 -129
rect -223 -163 -161 -129
rect -127 -163 -67 -129
rect -33 -163 31 -129
rect 65 -163 123 -129
rect 157 -163 223 -129
rect 257 -163 323 -129
rect 357 -163 383 -129
rect -377 -169 383 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +20 viadrn -20 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
