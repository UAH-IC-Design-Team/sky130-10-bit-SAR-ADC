magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< metal3 >>
rect -350 4432 349 4460
rect -350 78 265 4432
rect 329 78 349 4432
rect -350 50 349 78
rect -350 -78 349 -50
rect -350 -4432 265 -78
rect 329 -4432 349 -78
rect -350 -4460 349 -4432
<< via3 >>
rect 265 78 329 4432
rect 265 -4432 329 -78
<< mimcap >>
rect -250 4320 150 4360
rect -250 190 -210 4320
rect 110 190 150 4320
rect -250 150 150 190
rect -250 -190 150 -150
rect -250 -4320 -210 -190
rect 110 -4320 150 -190
rect -250 -4360 150 -4320
<< mimcapcontact >>
rect -210 190 110 4320
rect -210 -4320 110 -190
<< metal4 >>
rect -102 4321 2 4510
rect 218 4448 322 4510
rect 218 4432 345 4448
rect -211 4320 111 4321
rect -211 190 -210 4320
rect 110 190 111 4320
rect -211 189 111 190
rect -102 -189 2 189
rect 218 78 265 4432
rect 329 78 345 4432
rect 218 62 345 78
rect 218 -62 322 62
rect 218 -78 345 -62
rect -211 -190 111 -189
rect -211 -4320 -210 -190
rect 110 -4320 111 -190
rect -211 -4321 111 -4320
rect -102 -4510 2 -4321
rect 218 -4432 265 -78
rect 329 -4432 345 -78
rect 218 -4448 345 -4432
rect 218 -4510 322 -4448
<< properties >>
string FIXED_BBOX -350 50 250 4460
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
