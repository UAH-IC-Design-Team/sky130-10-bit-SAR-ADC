magic
tech sky130A
timestamp 1659111590
<< viali >>
rect 65 470 90 495
rect 345 475 375 500
rect 605 470 635 500
rect 170 440 195 465
rect 260 410 280 430
rect 25 385 50 402
rect 430 395 460 415
rect 520 410 540 430
<< metal1 >>
rect 125 520 160 570
rect 385 520 420 570
rect 645 520 685 570
rect 335 500 385 505
rect 55 495 205 500
rect 55 470 65 495
rect 90 470 205 495
rect 335 475 345 500
rect 375 475 385 500
rect 335 470 385 475
rect 595 500 645 505
rect 595 470 605 500
rect 635 470 645 500
rect 55 465 205 470
rect 595 465 645 470
rect 160 440 170 465
rect 195 440 205 465
rect 160 435 205 440
rect 250 434 550 455
rect 250 430 290 434
rect 250 410 260 430
rect 280 410 290 430
rect 510 430 550 434
rect 15 402 55 410
rect 250 405 290 410
rect 420 415 470 420
rect 15 385 25 402
rect 50 390 55 402
rect 420 395 430 415
rect 460 395 470 415
rect 510 410 520 430
rect 540 410 550 430
rect 510 405 550 410
rect 420 390 470 395
rect 50 385 470 390
rect 15 360 470 385
rect 125 250 160 300
rect 385 250 420 300
rect 645 250 685 300
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 684 0 1 274
box -19 -24 65 296
use sky130_fd_sc_hd__and2_0  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 159 0 1 274
box -19 -24 249 296
use sky130_fd_sc_hd__and2_0  x2
timestamp 1649977179
transform 1 0 419 0 1 274
box -19 -24 249 296
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 -11 0 1 274
box -19 -24 157 296
<< labels >>
rlabel metal1 140 570 140 570 5 VDD
port 1 s
rlabel metal1 135 250 135 250 1 VSS
port 2 n
rlabel metal1 140 360 140 360 1 S
port 3 n
rlabel metal1 365 435 365 435 1 IN
port 4 n
rlabel metal1 645 485 645 485 3 OUT_1
port 6 e
rlabel metal1 385 490 385 490 3 OUT_0
port 5 e
<< end >>
