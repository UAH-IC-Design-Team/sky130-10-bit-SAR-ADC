magic
tech sky130A
magscale 1 2
timestamp 1668294421
<< dnwell >>
rect 4600 400 6500 2300
<< nwell >>
rect 4520 2094 6580 2380
rect 4520 606 4806 2094
rect 6294 606 6580 2094
rect 4520 320 6580 606
<< nsubdiff >>
rect 4557 2323 6543 2343
rect 4557 2289 4637 2323
rect 6463 2289 6543 2323
rect 4557 2269 6543 2289
rect 4557 2263 4631 2269
rect 4557 437 4577 2263
rect 4611 437 4631 2263
rect 4557 431 4631 437
rect 6469 2263 6543 2269
rect 6469 437 6489 2263
rect 6523 437 6543 2263
rect 6469 431 6543 437
rect 4557 411 6543 431
rect 4557 377 4637 411
rect 6463 377 6543 411
rect 4557 357 6543 377
<< nsubdiffcont >>
rect 4637 2289 6463 2323
rect 4577 437 4611 2263
rect 6489 437 6523 2263
rect 4637 377 6463 411
<< locali >>
rect 4577 2289 4637 2323
rect 6463 2289 6523 2323
rect 4577 2263 4611 2289
rect 6489 2263 6523 2289
rect 5120 870 5950 880
rect 5120 790 5140 870
rect 5930 790 5950 870
rect 5120 780 5950 790
rect 4577 411 4611 437
rect 6489 411 6523 437
rect 4577 377 4637 411
rect 6463 377 6523 411
rect 5110 -830 5960 -820
rect 5110 -940 5130 -830
rect 5940 -940 5960 -830
rect 5110 -950 5960 -940
<< viali >>
rect 5140 790 5930 870
rect 5130 -940 5940 -830
<< metal1 >>
rect 5130 940 5950 1740
rect 5120 870 5950 880
rect 5120 790 5140 870
rect 5930 790 5950 870
rect 5120 -760 5950 790
rect 5110 -830 5960 -820
rect 5110 -940 5130 -830
rect 5940 -940 5960 -830
rect 5110 -950 5960 -940
use sky130_fd_pr__diode_pw2nd_05v5_EUY57X  D1
timestamp 1668293268
transform 1 0 5538 0 1 1338
box -538 -538 538 538
use sky130_fd_pr__diode_pw2nd_05v5_EUY57X  sky130_fd_pr__diode_pw2nd_05v5_EUY57X_0
timestamp 1668293268
transform 1 0 5538 0 1 -362
box -538 -538 538 538
<< labels >>
rlabel metal1 5130 940 5950 1740 1 VDD
port 1 n
rlabel metal1 5120 -760 5950 790 1 in
port 2 n
rlabel metal1 5110 -950 5960 -820 1 VSS
port 3 n
<< end >>
