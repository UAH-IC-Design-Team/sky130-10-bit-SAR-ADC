magic
tech sky130A
timestamp 1667684412
<< metal4 >>
rect 250 5200 310 5800
rect 590 5200 650 5800
rect 1050 5200 1110 5800
rect 1390 5200 1450 5800
rect 1850 5200 1910 5800
rect 2190 5200 2250 5800
rect 2650 5200 2710 5800
rect 2990 5200 3050 5800
rect 250 4400 310 5000
rect 590 4400 650 5000
rect 1050 4400 1110 5000
rect 1390 4400 1450 5000
rect 1850 4400 1910 5000
rect 2190 4400 2250 5000
rect 2650 4400 2710 5000
rect 2990 4400 3050 5000
rect 250 3600 310 4200
rect 590 3600 650 4200
rect 1050 3600 1110 4200
rect 1390 3600 1450 4200
rect 1850 3600 1910 4200
rect 2190 3600 2250 4200
rect 2650 3600 2710 4200
rect 2990 3600 3050 4200
rect 250 2800 310 3400
rect 590 2800 650 3400
rect 1050 2800 1110 3400
rect 1390 2800 1450 3400
rect 1850 2800 1910 3400
rect 2190 2800 2250 3400
rect 2650 2800 2710 3400
rect 2990 2800 3050 3400
rect 250 2000 310 2600
rect 590 2000 650 2600
rect 1050 2000 1110 2600
rect 1390 2000 1450 2600
rect 1850 2000 1910 2600
rect 2190 2000 2250 2600
rect 2650 2000 2710 2600
rect 2990 2000 3050 2600
rect 250 1200 310 1800
rect 590 1200 650 1800
rect 1050 1200 1110 1800
rect 1390 1200 1450 1800
rect 1850 1200 1910 1800
rect 2190 1200 2250 1800
rect 2650 1200 2710 1800
rect 2990 1200 3050 1800
rect 250 400 310 1000
rect 590 400 650 1000
rect 1050 400 1110 1000
rect 1390 400 1450 1000
rect 1850 400 1910 1000
rect 2190 400 2250 1000
rect 2650 400 2710 1000
rect 2990 400 3050 1000
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
array 0 3 800 0 7 800
timestamp 1667663783
transform 1 0 325 0 1 300
box -325 -300 325 300
<< end >>
