magic
tech sky130A
magscale 1 2
timestamp 1666552007
<< error_p >>
rect -269 246 -211 252
rect -77 246 -19 252
rect 115 246 173 252
rect 307 246 365 252
rect -269 212 -257 246
rect -77 212 -65 246
rect 115 212 127 246
rect 307 212 319 246
rect -269 206 -211 212
rect -77 206 -19 212
rect 115 206 173 212
rect 307 206 365 212
rect -365 -212 -307 -206
rect -173 -212 -115 -206
rect 19 -212 77 -206
rect 211 -212 269 -206
rect -365 -246 -353 -212
rect -173 -246 -161 -212
rect 19 -246 31 -212
rect 211 -246 223 -212
rect -365 -252 -307 -246
rect -173 -252 -115 -246
rect 19 -252 77 -246
rect 211 -252 269 -246
<< nwell >>
rect -353 227 449 265
rect -449 -227 449 227
rect -449 -265 353 -227
<< pmos >>
rect -351 -165 -321 165
rect -255 -165 -225 165
rect -159 -165 -129 165
rect -63 -165 -33 165
rect 33 -165 63 165
rect 129 -165 159 165
rect 225 -165 255 165
rect 321 -165 351 165
<< pdiff >>
rect -413 153 -351 165
rect -413 -153 -401 153
rect -367 -153 -351 153
rect -413 -165 -351 -153
rect -321 153 -255 165
rect -321 -153 -305 153
rect -271 -153 -255 153
rect -321 -165 -255 -153
rect -225 153 -159 165
rect -225 -153 -209 153
rect -175 -153 -159 153
rect -225 -165 -159 -153
rect -129 153 -63 165
rect -129 -153 -113 153
rect -79 -153 -63 153
rect -129 -165 -63 -153
rect -33 153 33 165
rect -33 -153 -17 153
rect 17 -153 33 153
rect -33 -165 33 -153
rect 63 153 129 165
rect 63 -153 79 153
rect 113 -153 129 153
rect 63 -165 129 -153
rect 159 153 225 165
rect 159 -153 175 153
rect 209 -153 225 153
rect 159 -165 225 -153
rect 255 153 321 165
rect 255 -153 271 153
rect 305 -153 321 153
rect 255 -165 321 -153
rect 351 153 413 165
rect 351 -153 367 153
rect 401 -153 413 153
rect 351 -165 413 -153
<< pdiffc >>
rect -401 -153 -367 153
rect -305 -153 -271 153
rect -209 -153 -175 153
rect -113 -153 -79 153
rect -17 -153 17 153
rect 79 -153 113 153
rect 175 -153 209 153
rect 271 -153 305 153
rect 367 -153 401 153
<< poly >>
rect -273 246 -207 262
rect -273 212 -257 246
rect -223 212 -207 246
rect -273 196 -207 212
rect -81 246 -15 262
rect -81 212 -65 246
rect -31 212 -15 246
rect -81 196 -15 212
rect 111 246 177 262
rect 111 212 127 246
rect 161 212 177 246
rect 111 196 177 212
rect 303 246 369 262
rect 303 212 319 246
rect 353 212 369 246
rect 303 196 369 212
rect -351 165 -321 191
rect -255 165 -225 196
rect -159 165 -129 191
rect -63 165 -33 196
rect 33 165 63 191
rect 129 165 159 196
rect 225 165 255 191
rect 321 165 351 196
rect -351 -196 -321 -165
rect -255 -191 -225 -165
rect -159 -196 -129 -165
rect -63 -191 -33 -165
rect 33 -196 63 -165
rect 129 -191 159 -165
rect 225 -196 255 -165
rect 321 -191 351 -165
rect -369 -212 -303 -196
rect -369 -246 -353 -212
rect -319 -246 -303 -212
rect -369 -262 -303 -246
rect -177 -212 -111 -196
rect -177 -246 -161 -212
rect -127 -246 -111 -212
rect -177 -262 -111 -246
rect 15 -212 81 -196
rect 15 -246 31 -212
rect 65 -246 81 -212
rect 15 -262 81 -246
rect 207 -212 273 -196
rect 207 -246 223 -212
rect 257 -246 273 -212
rect 207 -262 273 -246
<< polycont >>
rect -257 212 -223 246
rect -65 212 -31 246
rect 127 212 161 246
rect 319 212 353 246
rect -353 -246 -319 -212
rect -161 -246 -127 -212
rect 31 -246 65 -212
rect 223 -246 257 -212
<< locali >>
rect -273 212 -257 246
rect -223 212 -207 246
rect -81 212 -65 246
rect -31 212 -15 246
rect 111 212 127 246
rect 161 212 177 246
rect 303 212 319 246
rect 353 212 369 246
rect -401 153 -367 169
rect -401 -169 -367 -153
rect -305 153 -271 169
rect -305 -169 -271 -153
rect -209 153 -175 169
rect -209 -169 -175 -153
rect -113 153 -79 169
rect -113 -169 -79 -153
rect -17 153 17 169
rect -17 -169 17 -153
rect 79 153 113 169
rect 79 -169 113 -153
rect 175 153 209 169
rect 175 -169 209 -153
rect 271 153 305 169
rect 271 -169 305 -153
rect 367 153 401 169
rect 367 -169 401 -153
rect -369 -246 -353 -212
rect -319 -246 -303 -212
rect -177 -246 -161 -212
rect -127 -246 -111 -212
rect 15 -246 31 -212
rect 65 -246 81 -212
rect 207 -246 223 -212
rect 257 -246 273 -212
<< viali >>
rect -257 212 -223 246
rect -65 212 -31 246
rect 127 212 161 246
rect 319 212 353 246
rect -401 -153 -367 153
rect -305 -153 -271 153
rect -209 -153 -175 153
rect -113 -153 -79 153
rect -17 -153 17 153
rect 79 -153 113 153
rect 175 -153 209 153
rect 271 -153 305 153
rect 367 -153 401 153
rect -353 -246 -319 -212
rect -161 -246 -127 -212
rect 31 -246 65 -212
rect 223 -246 257 -212
<< metal1 >>
rect -269 246 -211 252
rect -269 212 -257 246
rect -223 212 -211 246
rect -269 206 -211 212
rect -77 246 -19 252
rect -77 212 -65 246
rect -31 212 -19 246
rect -77 206 -19 212
rect 115 246 173 252
rect 115 212 127 246
rect 161 212 173 246
rect 115 206 173 212
rect 307 246 365 252
rect 307 212 319 246
rect 353 212 365 246
rect 307 206 365 212
rect -407 153 -361 165
rect -407 -153 -401 153
rect -367 -153 -361 153
rect -407 -165 -361 -153
rect -311 153 -265 165
rect -311 -153 -305 153
rect -271 -153 -265 153
rect -311 -165 -265 -153
rect -215 153 -169 165
rect -215 -153 -209 153
rect -175 -153 -169 153
rect -215 -165 -169 -153
rect -119 153 -73 165
rect -119 -153 -113 153
rect -79 -153 -73 153
rect -119 -165 -73 -153
rect -23 153 23 165
rect -23 -153 -17 153
rect 17 -153 23 153
rect -23 -165 23 -153
rect 73 153 119 165
rect 73 -153 79 153
rect 113 -153 119 153
rect 73 -165 119 -153
rect 169 153 215 165
rect 169 -153 175 153
rect 209 -153 215 153
rect 169 -165 215 -153
rect 265 153 311 165
rect 265 -153 271 153
rect 305 -153 311 153
rect 265 -165 311 -153
rect 361 153 407 165
rect 361 -153 367 153
rect 401 -153 407 153
rect 361 -165 407 -153
rect -365 -212 -307 -206
rect -365 -246 -353 -212
rect -319 -246 -307 -212
rect -365 -252 -307 -246
rect -173 -212 -115 -206
rect -173 -246 -161 -212
rect -127 -246 -115 -212
rect -173 -252 -115 -246
rect 19 -212 77 -206
rect 19 -246 31 -212
rect 65 -246 77 -212
rect 19 -252 77 -246
rect 211 -212 269 -206
rect 211 -246 223 -212
rect 257 -246 269 -212
rect 211 -252 269 -246
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
