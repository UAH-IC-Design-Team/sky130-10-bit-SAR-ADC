magic
tech sky130A
magscale 1 2
timestamp 1665708526
<< error_s >>
rect 2712 7706 2770 7712
rect 2712 7672 2724 7706
rect 2712 7666 2770 7672
rect 2712 7598 2770 7604
rect 2712 7564 2724 7598
rect 2712 7558 2770 7564
rect 2712 7140 2770 7146
rect 2712 7106 2724 7140
rect 2712 7100 2770 7106
rect 2712 7032 2770 7038
rect 2712 6998 2724 7032
rect 2712 6992 2770 6998
rect 2566 6831 2600 6849
rect 2343 6693 2401 6699
rect 2343 6659 2355 6693
rect 2343 6653 2401 6659
rect 2343 6401 2401 6407
rect 2343 6367 2355 6401
rect 2343 6361 2401 6367
rect 2343 6293 2401 6299
rect 2343 6259 2355 6293
rect 2343 6253 2401 6259
rect 2343 6001 2401 6007
rect 2343 5967 2355 6001
rect 2343 5961 2401 5967
rect 2343 5893 2401 5899
rect 2343 5859 2355 5893
rect 2343 5853 2401 5859
rect 2343 5601 2401 5607
rect 2343 5567 2355 5601
rect 2343 5561 2401 5567
rect 2343 5493 2401 5499
rect 2343 5459 2355 5493
rect 2343 5453 2401 5459
rect 2343 5201 2401 5207
rect 2343 5167 2355 5201
rect 2343 5161 2401 5167
rect 2343 5093 2401 5099
rect 2343 5059 2355 5093
rect 2343 5053 2401 5059
rect 2197 5012 2231 5030
rect 1974 4874 2032 4880
rect 1974 4840 1986 4874
rect 1974 4834 2032 4840
rect 1974 4416 2032 4422
rect 1974 4382 1986 4416
rect 1974 4376 2032 4382
rect 1974 4308 2032 4314
rect 1974 4274 1986 4308
rect 1974 4268 2032 4274
rect 1974 3850 2032 3856
rect 1974 3816 1986 3850
rect 1974 3810 2032 3816
rect 1828 3737 1862 3755
rect 1605 3599 1663 3605
rect 1605 3565 1617 3599
rect 1605 3559 1663 3565
rect 1605 3307 1663 3313
rect 1605 3273 1617 3307
rect 1605 3267 1663 3273
rect 1605 3199 1663 3205
rect 1605 3165 1617 3199
rect 1605 3159 1663 3165
rect 1605 2907 1663 2913
rect 1605 2873 1617 2907
rect 1459 2854 1493 2872
rect 1605 2867 1663 2873
rect 1236 2716 1294 2722
rect 1236 2682 1248 2716
rect 1236 2676 1294 2682
rect 1090 2243 1124 2261
rect 867 2105 925 2111
rect 867 2071 879 2105
rect 867 2065 925 2071
rect 867 1813 925 1819
rect 867 1779 879 1813
rect 867 1773 925 1779
rect 867 1705 925 1711
rect 867 1671 879 1705
rect 867 1665 925 1671
rect 867 1413 925 1419
rect 867 1379 879 1413
rect 867 1373 925 1379
rect 867 1305 925 1311
rect 721 1262 755 1280
rect 867 1271 879 1305
rect 867 1265 925 1271
rect 352 1149 386 1167
rect 129 1011 187 1017
rect 129 977 141 1011
rect 129 971 187 977
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1149
rect 498 1124 556 1130
rect 498 1090 510 1124
rect 498 1084 556 1090
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 685 530 755 1262
rect 867 1013 925 1019
rect 867 979 879 1013
rect 867 973 925 979
rect 867 905 925 911
rect 867 871 879 905
rect 867 865 925 871
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1054 477 1124 2243
rect 1236 2258 1294 2264
rect 1236 2224 1248 2258
rect 1236 2218 1294 2224
rect 1236 2150 1294 2156
rect 1236 2116 1248 2150
rect 1236 2110 1294 2116
rect 1236 1692 1294 1698
rect 1236 1658 1248 1692
rect 1236 1652 1294 1658
rect 1236 1584 1294 1590
rect 1236 1550 1248 1584
rect 1236 1544 1294 1550
rect 1236 1126 1294 1132
rect 1236 1092 1248 1126
rect 1236 1086 1294 1092
rect 1236 1018 1294 1024
rect 1236 984 1248 1018
rect 1236 978 1294 984
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1054 441 1107 477
rect 1423 424 1493 2854
rect 1605 2799 1663 2805
rect 1605 2765 1617 2799
rect 1605 2759 1663 2765
rect 1605 2507 1663 2513
rect 1605 2473 1617 2507
rect 1605 2467 1663 2473
rect 1605 2399 1663 2405
rect 1605 2365 1617 2399
rect 1605 2359 1663 2365
rect 1605 2107 1663 2113
rect 1605 2073 1617 2107
rect 1605 2067 1663 2073
rect 1605 1999 1663 2005
rect 1605 1965 1617 1999
rect 1605 1959 1663 1965
rect 1605 1707 1663 1713
rect 1605 1673 1617 1707
rect 1605 1667 1663 1673
rect 1605 1599 1663 1605
rect 1605 1565 1617 1599
rect 1605 1559 1663 1565
rect 1605 1307 1663 1313
rect 1605 1273 1617 1307
rect 1605 1267 1663 1273
rect 1605 1199 1663 1205
rect 1605 1165 1617 1199
rect 1605 1159 1663 1165
rect 1605 907 1663 913
rect 1605 873 1617 907
rect 1605 867 1663 873
rect 1605 799 1663 805
rect 1605 765 1617 799
rect 1605 759 1663 765
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1792 371 1862 3737
rect 1974 3742 2032 3748
rect 1974 3708 1986 3742
rect 1974 3702 2032 3708
rect 1974 3284 2032 3290
rect 1974 3250 1986 3284
rect 1974 3244 2032 3250
rect 1974 3176 2032 3182
rect 1974 3142 1986 3176
rect 1974 3136 2032 3142
rect 1974 2718 2032 2724
rect 1974 2684 1986 2718
rect 1974 2678 2032 2684
rect 1974 2610 2032 2616
rect 1974 2576 1986 2610
rect 1974 2570 2032 2576
rect 1974 2152 2032 2158
rect 1974 2118 1986 2152
rect 1974 2112 2032 2118
rect 1974 2044 2032 2050
rect 1974 2010 1986 2044
rect 1974 2004 2032 2010
rect 1974 1586 2032 1592
rect 1974 1552 1986 1586
rect 1974 1546 2032 1552
rect 1974 1478 2032 1484
rect 1974 1444 1986 1478
rect 1974 1438 2032 1444
rect 1974 1020 2032 1026
rect 1974 986 1986 1020
rect 1974 980 2032 986
rect 1974 912 2032 918
rect 1974 878 1986 912
rect 1974 872 2032 878
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
rect 2161 318 2231 5012
rect 2343 4801 2401 4807
rect 2343 4767 2355 4801
rect 2343 4761 2401 4767
rect 2343 4693 2401 4699
rect 2343 4659 2355 4693
rect 2343 4653 2401 4659
rect 2343 4401 2401 4407
rect 2343 4367 2355 4401
rect 2343 4361 2401 4367
rect 2343 4293 2401 4299
rect 2343 4259 2355 4293
rect 2343 4253 2401 4259
rect 2343 4001 2401 4007
rect 2343 3967 2355 4001
rect 2343 3961 2401 3967
rect 2343 3893 2401 3899
rect 2343 3859 2355 3893
rect 2343 3853 2401 3859
rect 2343 3601 2401 3607
rect 2343 3567 2355 3601
rect 2343 3561 2401 3567
rect 2343 3493 2401 3499
rect 2343 3459 2355 3493
rect 2343 3453 2401 3459
rect 2343 3201 2401 3207
rect 2343 3167 2355 3201
rect 2343 3161 2401 3167
rect 2343 3093 2401 3099
rect 2343 3059 2355 3093
rect 2343 3053 2401 3059
rect 2343 2801 2401 2807
rect 2343 2767 2355 2801
rect 2343 2761 2401 2767
rect 2343 2693 2401 2699
rect 2343 2659 2355 2693
rect 2343 2653 2401 2659
rect 2343 2401 2401 2407
rect 2343 2367 2355 2401
rect 2343 2361 2401 2367
rect 2343 2293 2401 2299
rect 2343 2259 2355 2293
rect 2343 2253 2401 2259
rect 2343 2001 2401 2007
rect 2343 1967 2355 2001
rect 2343 1961 2401 1967
rect 2343 1893 2401 1899
rect 2343 1859 2355 1893
rect 2343 1853 2401 1859
rect 2343 1601 2401 1607
rect 2343 1567 2355 1601
rect 2343 1561 2401 1567
rect 2343 1493 2401 1499
rect 2343 1459 2355 1493
rect 2343 1453 2401 1459
rect 2343 1201 2401 1207
rect 2343 1167 2355 1201
rect 2343 1161 2401 1167
rect 2343 1093 2401 1099
rect 2343 1059 2355 1093
rect 2343 1053 2401 1059
rect 2343 801 2401 807
rect 2343 767 2355 801
rect 2343 761 2401 767
rect 2343 693 2401 699
rect 2343 659 2355 693
rect 2343 653 2401 659
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2161 282 2214 318
rect 2530 265 2600 6831
rect 2712 6574 2770 6580
rect 2712 6540 2724 6574
rect 2712 6534 2770 6540
rect 2712 6466 2770 6472
rect 2712 6432 2724 6466
rect 2712 6426 2770 6432
rect 2712 6008 2770 6014
rect 2712 5974 2724 6008
rect 2712 5968 2770 5974
rect 2712 5900 2770 5906
rect 2712 5866 2724 5900
rect 2712 5860 2770 5866
rect 2712 5442 2770 5448
rect 2712 5408 2724 5442
rect 2712 5402 2770 5408
rect 2712 5334 2770 5340
rect 2712 5300 2724 5334
rect 2712 5294 2770 5300
rect 2712 4876 2770 4882
rect 2712 4842 2724 4876
rect 2712 4836 2770 4842
rect 2712 4768 2770 4774
rect 2712 4734 2724 4768
rect 2712 4728 2770 4734
rect 2712 4310 2770 4316
rect 2712 4276 2724 4310
rect 2712 4270 2770 4276
rect 2712 4202 2770 4208
rect 2712 4168 2724 4202
rect 2712 4162 2770 4168
rect 2712 3744 2770 3750
rect 2712 3710 2724 3744
rect 2712 3704 2770 3710
rect 2712 3636 2770 3642
rect 2712 3602 2724 3636
rect 2712 3596 2770 3602
rect 2712 3178 2770 3184
rect 2712 3144 2724 3178
rect 2712 3138 2770 3144
rect 2712 3070 2770 3076
rect 2712 3036 2724 3070
rect 2712 3030 2770 3036
rect 2712 2612 2770 2618
rect 2712 2578 2724 2612
rect 2712 2572 2770 2578
rect 2712 2504 2770 2510
rect 2712 2470 2724 2504
rect 2712 2464 2770 2470
rect 2712 2046 2770 2052
rect 2712 2012 2724 2046
rect 2712 2006 2770 2012
rect 2712 1938 2770 1944
rect 2712 1904 2724 1938
rect 2712 1898 2770 1904
rect 2712 1480 2770 1486
rect 2712 1446 2724 1480
rect 2712 1440 2770 1446
rect 2712 1372 2770 1378
rect 2712 1338 2724 1372
rect 2712 1332 2770 1338
rect 2712 914 2770 920
rect 2712 880 2724 914
rect 2712 874 2770 880
rect 2712 806 2770 812
rect 2712 772 2724 806
rect 2712 766 2770 772
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2530 229 2583 265
<< metal4 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_77T378  XM1
timestamp 1665708526
transform 1 0 158 0 1 848
box -211 -301 211 301
use sky130_fd_pr__pfet_01v8_XJF7MR  XM2
timestamp 1665708526
transform 1 0 527 0 1 878
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_YBY378  XM3
timestamp 1665708526
transform 1 0 896 0 1 1342
box -211 -901 211 901
use sky130_fd_pr__pfet_01v8_KJFHF3  XM4
timestamp 1665708526
transform 1 0 1265 0 1 1621
box -211 -1233 211 1233
use sky130_fd_pr__nfet_01v8_CCZD88  XM5
timestamp 1665708526
transform 1 0 1634 0 1 2036
box -211 -1701 211 1701
use sky130_fd_pr__pfet_01v8_MJF9NY  XM6
timestamp 1665708526
transform 1 0 2003 0 1 2647
box -211 -2365 211 2365
use sky130_fd_pr__nfet_01v8_UDP43T  XM7
timestamp 1665708526
transform 1 0 2372 0 1 3530
box -211 -3301 211 3301
use sky130_fd_pr__pfet_01v8_UNNRDR  XM8
timestamp 1665708526
transform 1 0 2741 0 1 4805
box -211 -4629 211 4629
<< labels >>
flabel metal4 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal4 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal4 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal4 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
