magic
tech sky130A
magscale 1 2
timestamp 1668016263
<< nwell >>
rect -300 1100 1690 2810
<< psubdiff >>
rect -140 790 -30 814
rect -140 656 -30 680
rect -14 540 10 600
rect 180 540 204 600
rect 300 460 370 484
rect 300 316 370 340
rect 396 120 420 190
rect 590 120 614 190
rect 800 20 870 44
rect 800 -144 870 -120
rect 916 -650 940 -580
rect 1150 -650 1174 -580
<< nsubdiff >>
rect 820 2620 850 2690
rect 940 2620 970 2690
rect 820 2340 850 2410
rect 940 2340 970 2410
rect 820 2090 850 2160
rect 940 2090 970 2160
rect 320 1830 350 1900
rect 440 1830 470 1900
rect 320 1680 350 1750
rect 440 1680 470 1750
rect -30 1480 0 1550
rect 100 1480 130 1550
rect -30 1350 0 1420
rect 100 1350 130 1420
<< psubdiffcont >>
rect -140 680 -30 790
rect 10 540 180 600
rect 300 340 370 460
rect 420 120 590 190
rect 800 -120 870 20
rect 940 -650 1150 -580
<< nsubdiffcont >>
rect 850 2620 940 2690
rect 850 2340 940 2410
rect 850 2090 940 2160
rect 350 1830 440 1900
rect 350 1680 440 1750
rect 0 1480 100 1550
rect 0 1350 100 1420
<< locali >>
rect 830 2620 850 2690
rect 940 2620 960 2690
rect 830 2340 850 2410
rect 940 2340 960 2410
rect 830 2090 850 2160
rect 940 2090 960 2160
rect 330 1830 350 1900
rect 440 1830 460 1900
rect 330 1680 350 1750
rect 440 1680 460 1750
rect -20 1480 0 1550
rect 100 1480 120 1550
rect -20 1350 0 1420
rect 100 1350 120 1420
rect -140 790 -30 806
rect -140 670 -130 680
rect -40 670 -30 680
rect -140 664 -30 670
rect -6 540 10 600
rect 180 540 196 600
rect 300 460 370 476
rect 300 324 370 340
rect 404 120 420 190
rect 590 120 606 190
rect 800 20 870 36
rect 800 -136 870 -120
rect 924 -650 940 -580
rect 1150 -650 1166 -580
<< viali >>
rect 850 2620 940 2690
rect 850 2340 940 2410
rect 850 2090 940 2160
rect 350 1830 440 1900
rect 350 1680 440 1750
rect 0 1480 100 1550
rect 0 1350 100 1420
rect -130 680 -40 790
rect -130 670 -40 680
rect 20 550 170 590
rect 310 350 360 450
rect 430 130 580 180
rect 810 -110 860 10
rect 950 -640 1140 -590
<< metal1 >>
rect 840 2740 1450 2810
rect 840 2690 950 2740
rect 840 2620 850 2690
rect 940 2620 950 2690
rect 840 2410 950 2620
rect 840 2340 850 2410
rect 940 2340 950 2410
rect 840 2160 950 2340
rect 840 2090 850 2160
rect 940 2090 950 2160
rect 840 2060 950 2090
rect 340 1990 950 2060
rect 340 1900 450 1990
rect 340 1830 350 1900
rect 440 1830 450 1900
rect 340 1750 450 1830
rect 340 1680 350 1750
rect 440 1680 450 1750
rect 340 1660 450 1680
rect -10 1590 450 1660
rect -10 1550 110 1590
rect -10 1480 0 1550
rect 100 1480 110 1550
rect -10 1420 110 1480
rect -10 1350 0 1420
rect 100 1350 110 1420
rect -290 920 -240 1250
rect -10 1230 110 1350
rect -190 1100 -40 1180
rect 230 1100 280 1540
rect 340 1240 450 1590
rect 530 1100 640 1570
rect 730 1100 780 1930
rect 840 1240 950 1990
rect 1020 1100 1130 1950
rect 1230 1100 1280 2690
rect 1340 1240 1450 2740
rect 1520 1100 1730 2730
rect -190 1060 280 1100
rect -190 980 -40 1060
rect -140 790 -30 930
rect -140 670 -130 790
rect -40 670 -30 790
rect -140 600 -30 670
rect 230 630 280 1060
rect 430 1060 780 1100
rect 310 600 370 930
rect -140 590 370 600
rect 430 590 480 1060
rect -140 550 20 590
rect 170 550 370 590
rect -140 540 370 550
rect 300 450 370 540
rect 300 350 310 450
rect 360 350 370 450
rect 300 190 370 350
rect 730 230 780 1060
rect 930 1060 1280 1100
rect 810 190 870 930
rect 930 200 990 1060
rect 300 180 870 190
rect 300 130 430 180
rect 580 130 870 180
rect 300 120 870 130
rect 800 10 870 120
rect 800 -110 810 10
rect 860 -110 870 10
rect 800 -580 870 -110
rect 1230 -540 1280 1060
rect 1430 1090 1730 1100
rect 1430 1030 1650 1090
rect 1310 -580 1370 920
rect 1430 -570 1630 1030
rect 800 -590 1370 -580
rect 800 -640 950 -590
rect 1140 -640 1370 -590
rect 800 -650 1370 -640
use sky130_fd_pr__pfet_01v8_BBAHKR  XM4
timestamp 1666553317
transform 0 1 485 -1 0 1357
box -263 -265 257 205
use sky130_fd_pr__nfet_01v8_HRFJZU  XM5
timestamp 1666552870
transform 0 1 899 -1 0 613
box -413 -179 413 121
use sky130_fd_pr__pfet_01v8_BBSRKR  XM6
timestamp 1666553528
transform 0 1 985 -1 0 1549
box -451 -265 449 205
use sky130_fd_pr__nfet_01v8_29RM5N  XM7
timestamp 1667868113
transform 0 1 1399 -1 0 227
box -797 -179 797 121
use sky130_fd_pr__pfet_01v8_2FR7QD  XM8
timestamp 1666553750
transform 0 1 1485 -1 0 1933
box -837 -265 833 205
use sky130_fd_pr__nfet_01v8_5EDJZL  sky130_fd_pr__nfet_01v8_5EDJZL_0
timestamp 1666555252
transform 0 1 399 -1 0 811
box -221 -179 221 121
use sky130_fd_pr__nfet_01v8_9CGS2F  sky130_fd_pr__nfet_01v8_9CGS2F_0
timestamp 1666651042
transform 0 1 -152 -1 0 953
box -73 -148 73 148
use sky130_fd_pr__pfet_01v8_46WN3R  sky130_fd_pr__pfet_01v8_46WN3R_0
timestamp 1666487809
transform 0 1 -71 1 0 1209
box -109 -229 109 263
<< end >>
