magic
tech sky130A
magscale 1 2
timestamp 1665780148
<< error_p >>
rect -29 375 29 381
rect -29 341 -17 375
rect -29 335 29 341
<< nwell >>
rect -109 -428 109 394
<< pmos >>
rect -15 -366 15 294
<< pdiff >>
rect -73 282 -15 294
rect -73 -354 -61 282
rect -27 -354 -15 282
rect -73 -366 -15 -354
rect 15 282 73 294
rect 15 -354 27 282
rect 61 -354 73 282
rect 15 -366 73 -354
<< pdiffc >>
rect -61 -354 -27 282
rect 27 -354 61 282
<< poly >>
rect -33 375 33 391
rect -33 341 -17 375
rect 17 341 33 375
rect -33 325 33 341
rect -15 294 15 325
rect -15 -392 15 -366
<< polycont >>
rect -17 341 17 375
<< locali >>
rect -33 341 -17 375
rect 17 341 33 375
rect -61 282 -27 298
rect -61 -370 -27 -354
rect 27 282 61 298
rect 27 -370 61 -354
<< viali >>
rect -17 341 17 375
rect -61 11 -27 265
rect 27 -354 61 282
<< metal1 >>
rect -29 375 29 381
rect -29 341 -17 375
rect 17 341 29 375
rect -29 335 29 341
rect 21 282 67 294
rect -67 265 -21 277
rect -67 11 -61 265
rect -27 11 -21 265
rect -67 -1 -21 11
rect 21 -354 27 282
rect 61 -354 67 282
rect 21 -366 67 -354
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.3 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
