magic
tech sky130A
magscale 1 2
timestamp 1668018737
<< nwell >>
rect -300 910 730 1240
rect -300 900 240 910
<< psubdiff >>
rect 70 780 130 804
rect 70 656 130 680
<< nsubdiff >>
rect -200 1190 -100 1200
rect -200 1150 -170 1190
rect -130 1150 -100 1190
rect -200 1140 -100 1150
rect -10 1190 90 1200
rect -10 1150 20 1190
rect 60 1150 90 1190
rect -10 1140 90 1150
<< psubdiffcont >>
rect 70 680 130 780
<< nsubdiffcont >>
rect -170 1150 -130 1190
rect 20 1150 60 1190
<< locali >>
rect -190 1190 -110 1200
rect -190 1150 -170 1190
rect -130 1150 -110 1190
rect -190 1140 -110 1150
rect 0 1190 80 1200
rect 0 1150 20 1190
rect 60 1150 80 1190
rect 0 1140 80 1150
rect 70 780 130 796
rect 70 664 130 680
<< viali >>
rect -170 1150 -130 1190
rect 20 1150 60 1190
rect 80 690 120 770
<< metal1 >>
rect -190 1190 -110 1200
rect -190 1150 -170 1190
rect -130 1150 -110 1190
rect -190 1110 -110 1150
rect 0 1190 380 1210
rect 0 1150 20 1190
rect 60 1170 380 1190
rect 60 1150 80 1170
rect 0 1110 80 1150
rect -200 1070 130 1110
rect -300 720 -240 1040
rect -200 910 -40 980
rect 200 910 260 1140
rect 330 1040 380 1170
rect -200 850 260 910
rect -200 780 -40 850
rect 70 770 130 790
rect 70 720 80 770
rect 50 690 80 720
rect 120 720 130 770
rect 200 720 260 850
rect 480 780 640 1180
rect 120 690 150 720
rect -200 650 650 690
use sky130_fd_pr__nfet_01v8_9CME3F  XM1
timestamp 1666651042
transform 0 -1 -152 1 0 753
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_Z2KCLS  XM3
timestamp 1665882771
transform 0 -1 439 1 0 753
box -73 -239 73 239
use sky130_fd_pr__pfet_01v8_5AWN3K  sky130_fd_pr__pfet_01v8_5AWN3K_0
timestamp 1665779562
transform 0 -1 -71 1 0 1009
box -109 -263 109 229
use sky130_fd_pr__pfet_01v8_S6MTYS  sky130_fd_pr__pfet_01v8_S6MTYS_0
timestamp 1666374753
transform 0 -1 465 1 0 1061
box -161 -265 177 265
<< labels >>
rlabel metal1 -200 1070 130 1110 1 VDD
port 1 n
rlabel metal1 -300 720 -240 1040 1 Vin
port 2 n
rlabel metal1 480 780 620 1180 1 Vout
port 3 n
rlabel metal1 -200 650 650 690 1 VSS
port 4 n
<< end >>
