magic
tech sky130A
magscale 1 2
timestamp 1665159686
<< metal3 >>
rect -350 36002 349 36030
rect -350 31648 265 36002
rect 329 31648 349 36002
rect -350 31620 349 31648
rect -350 31492 349 31520
rect -350 27138 265 31492
rect 329 27138 349 31492
rect -350 27110 349 27138
rect -350 26982 349 27010
rect -350 22628 265 26982
rect 329 22628 349 26982
rect -350 22600 349 22628
rect -350 22472 349 22500
rect -350 18118 265 22472
rect 329 18118 349 22472
rect -350 18090 349 18118
rect -350 17962 349 17990
rect -350 13608 265 17962
rect 329 13608 349 17962
rect -350 13580 349 13608
rect -350 13452 349 13480
rect -350 9098 265 13452
rect 329 9098 349 13452
rect -350 9070 349 9098
rect -350 8942 349 8970
rect -350 4588 265 8942
rect 329 4588 349 8942
rect -350 4560 349 4588
rect -350 4432 349 4460
rect -350 78 265 4432
rect 329 78 349 4432
rect -350 50 349 78
rect -350 -78 349 -50
rect -350 -4432 265 -78
rect 329 -4432 349 -78
rect -350 -4460 349 -4432
rect -350 -4588 349 -4560
rect -350 -8942 265 -4588
rect 329 -8942 349 -4588
rect -350 -8970 349 -8942
rect -350 -9098 349 -9070
rect -350 -13452 265 -9098
rect 329 -13452 349 -9098
rect -350 -13480 349 -13452
rect -350 -13608 349 -13580
rect -350 -17962 265 -13608
rect 329 -17962 349 -13608
rect -350 -17990 349 -17962
rect -350 -18118 349 -18090
rect -350 -22472 265 -18118
rect 329 -22472 349 -18118
rect -350 -22500 349 -22472
rect -350 -22628 349 -22600
rect -350 -26982 265 -22628
rect 329 -26982 349 -22628
rect -350 -27010 349 -26982
rect -350 -27138 349 -27110
rect -350 -31492 265 -27138
rect 329 -31492 349 -27138
rect -350 -31520 349 -31492
rect -350 -31648 349 -31620
rect -350 -36002 265 -31648
rect 329 -36002 349 -31648
rect -350 -36030 349 -36002
<< via3 >>
rect 265 31648 329 36002
rect 265 27138 329 31492
rect 265 22628 329 26982
rect 265 18118 329 22472
rect 265 13608 329 17962
rect 265 9098 329 13452
rect 265 4588 329 8942
rect 265 78 329 4432
rect 265 -4432 329 -78
rect 265 -8942 329 -4588
rect 265 -13452 329 -9098
rect 265 -17962 329 -13608
rect 265 -22472 329 -18118
rect 265 -26982 329 -22628
rect 265 -31492 329 -27138
rect 265 -36002 329 -31648
<< mimcap >>
rect -250 35890 150 35930
rect -250 31760 -210 35890
rect 110 31760 150 35890
rect -250 31720 150 31760
rect -250 31380 150 31420
rect -250 27250 -210 31380
rect 110 27250 150 31380
rect -250 27210 150 27250
rect -250 26870 150 26910
rect -250 22740 -210 26870
rect 110 22740 150 26870
rect -250 22700 150 22740
rect -250 22360 150 22400
rect -250 18230 -210 22360
rect 110 18230 150 22360
rect -250 18190 150 18230
rect -250 17850 150 17890
rect -250 13720 -210 17850
rect 110 13720 150 17850
rect -250 13680 150 13720
rect -250 13340 150 13380
rect -250 9210 -210 13340
rect 110 9210 150 13340
rect -250 9170 150 9210
rect -250 8830 150 8870
rect -250 4700 -210 8830
rect 110 4700 150 8830
rect -250 4660 150 4700
rect -250 4320 150 4360
rect -250 190 -210 4320
rect 110 190 150 4320
rect -250 150 150 190
rect -250 -190 150 -150
rect -250 -4320 -210 -190
rect 110 -4320 150 -190
rect -250 -4360 150 -4320
rect -250 -4700 150 -4660
rect -250 -8830 -210 -4700
rect 110 -8830 150 -4700
rect -250 -8870 150 -8830
rect -250 -9210 150 -9170
rect -250 -13340 -210 -9210
rect 110 -13340 150 -9210
rect -250 -13380 150 -13340
rect -250 -13720 150 -13680
rect -250 -17850 -210 -13720
rect 110 -17850 150 -13720
rect -250 -17890 150 -17850
rect -250 -18230 150 -18190
rect -250 -22360 -210 -18230
rect 110 -22360 150 -18230
rect -250 -22400 150 -22360
rect -250 -22740 150 -22700
rect -250 -26870 -210 -22740
rect 110 -26870 150 -22740
rect -250 -26910 150 -26870
rect -250 -27250 150 -27210
rect -250 -31380 -210 -27250
rect 110 -31380 150 -27250
rect -250 -31420 150 -31380
rect -250 -31760 150 -31720
rect -250 -35890 -210 -31760
rect 110 -35890 150 -31760
rect -250 -35930 150 -35890
<< mimcapcontact >>
rect -210 31760 110 35890
rect -210 27250 110 31380
rect -210 22740 110 26870
rect -210 18230 110 22360
rect -210 13720 110 17850
rect -210 9210 110 13340
rect -210 4700 110 8830
rect -210 190 110 4320
rect -210 -4320 110 -190
rect -210 -8830 110 -4700
rect -210 -13340 110 -9210
rect -210 -17850 110 -13720
rect -210 -22360 110 -18230
rect -210 -26870 110 -22740
rect -210 -31380 110 -27250
rect -210 -35890 110 -31760
<< metal4 >>
rect -102 35891 2 36080
rect 218 36018 322 36080
rect 218 36002 345 36018
rect -211 35890 111 35891
rect -211 31760 -210 35890
rect 110 31760 111 35890
rect -211 31759 111 31760
rect -102 31381 2 31759
rect 218 31648 265 36002
rect 329 31648 345 36002
rect 218 31632 345 31648
rect 218 31508 322 31632
rect 218 31492 345 31508
rect -211 31380 111 31381
rect -211 27250 -210 31380
rect 110 27250 111 31380
rect -211 27249 111 27250
rect -102 26871 2 27249
rect 218 27138 265 31492
rect 329 27138 345 31492
rect 218 27122 345 27138
rect 218 26998 322 27122
rect 218 26982 345 26998
rect -211 26870 111 26871
rect -211 22740 -210 26870
rect 110 22740 111 26870
rect -211 22739 111 22740
rect -102 22361 2 22739
rect 218 22628 265 26982
rect 329 22628 345 26982
rect 218 22612 345 22628
rect 218 22488 322 22612
rect 218 22472 345 22488
rect -211 22360 111 22361
rect -211 18230 -210 22360
rect 110 18230 111 22360
rect -211 18229 111 18230
rect -102 17851 2 18229
rect 218 18118 265 22472
rect 329 18118 345 22472
rect 218 18102 345 18118
rect 218 17978 322 18102
rect 218 17962 345 17978
rect -211 17850 111 17851
rect -211 13720 -210 17850
rect 110 13720 111 17850
rect -211 13719 111 13720
rect -102 13341 2 13719
rect 218 13608 265 17962
rect 329 13608 345 17962
rect 218 13592 345 13608
rect 218 13468 322 13592
rect 218 13452 345 13468
rect -211 13340 111 13341
rect -211 9210 -210 13340
rect 110 9210 111 13340
rect -211 9209 111 9210
rect -102 8831 2 9209
rect 218 9098 265 13452
rect 329 9098 345 13452
rect 218 9082 345 9098
rect 218 8958 322 9082
rect 218 8942 345 8958
rect -211 8830 111 8831
rect -211 4700 -210 8830
rect 110 4700 111 8830
rect -211 4699 111 4700
rect -102 4321 2 4699
rect 218 4588 265 8942
rect 329 4588 345 8942
rect 218 4572 345 4588
rect 218 4448 322 4572
rect 218 4432 345 4448
rect -211 4320 111 4321
rect -211 190 -210 4320
rect 110 190 111 4320
rect -211 189 111 190
rect -102 -189 2 189
rect 218 78 265 4432
rect 329 78 345 4432
rect 218 62 345 78
rect 218 -62 322 62
rect 218 -78 345 -62
rect -211 -190 111 -189
rect -211 -4320 -210 -190
rect 110 -4320 111 -190
rect -211 -4321 111 -4320
rect -102 -4699 2 -4321
rect 218 -4432 265 -78
rect 329 -4432 345 -78
rect 218 -4448 345 -4432
rect 218 -4572 322 -4448
rect 218 -4588 345 -4572
rect -211 -4700 111 -4699
rect -211 -8830 -210 -4700
rect 110 -8830 111 -4700
rect -211 -8831 111 -8830
rect -102 -9209 2 -8831
rect 218 -8942 265 -4588
rect 329 -8942 345 -4588
rect 218 -8958 345 -8942
rect 218 -9082 322 -8958
rect 218 -9098 345 -9082
rect -211 -9210 111 -9209
rect -211 -13340 -210 -9210
rect 110 -13340 111 -9210
rect -211 -13341 111 -13340
rect -102 -13719 2 -13341
rect 218 -13452 265 -9098
rect 329 -13452 345 -9098
rect 218 -13468 345 -13452
rect 218 -13592 322 -13468
rect 218 -13608 345 -13592
rect -211 -13720 111 -13719
rect -211 -17850 -210 -13720
rect 110 -17850 111 -13720
rect -211 -17851 111 -17850
rect -102 -18229 2 -17851
rect 218 -17962 265 -13608
rect 329 -17962 345 -13608
rect 218 -17978 345 -17962
rect 218 -18102 322 -17978
rect 218 -18118 345 -18102
rect -211 -18230 111 -18229
rect -211 -22360 -210 -18230
rect 110 -22360 111 -18230
rect -211 -22361 111 -22360
rect -102 -22739 2 -22361
rect 218 -22472 265 -18118
rect 329 -22472 345 -18118
rect 218 -22488 345 -22472
rect 218 -22612 322 -22488
rect 218 -22628 345 -22612
rect -211 -22740 111 -22739
rect -211 -26870 -210 -22740
rect 110 -26870 111 -22740
rect -211 -26871 111 -26870
rect -102 -27249 2 -26871
rect 218 -26982 265 -22628
rect 329 -26982 345 -22628
rect 218 -26998 345 -26982
rect 218 -27122 322 -26998
rect 218 -27138 345 -27122
rect -211 -27250 111 -27249
rect -211 -31380 -210 -27250
rect 110 -31380 111 -27250
rect -211 -31381 111 -31380
rect -102 -31759 2 -31381
rect 218 -31492 265 -27138
rect 329 -31492 345 -27138
rect 218 -31508 345 -31492
rect 218 -31632 322 -31508
rect 218 -31648 345 -31632
rect -211 -31760 111 -31759
rect -211 -35890 -210 -31760
rect 110 -35890 111 -31760
rect -211 -35891 111 -35890
rect -102 -36080 2 -35891
rect 218 -36002 265 -31648
rect 329 -36002 345 -31648
rect 218 -36018 345 -36002
rect 218 -36080 322 -36018
<< properties >>
string FIXED_BBOX -350 31620 250 36030
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.97 carea 2.00 cperi 0.19 nx 1 ny 16 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
