* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
** sch_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/tests/pulse_generator/pulse_generator_test.sch
**.subckt pulse_generator_test
**** begin user architecture code
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
**** end user architecture code
**.ends
* expanding   symbol:  src/pulse_generator/pulse_generator.sym # of pins=5
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/pulse_generator/pulse_generator.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/pulse_generator/pulse_generator.sch
.subckt pulse_generator a_clk a_pulse a_VDD a_VSS a_RST_PLS
*.ipin clk
*.ipin RST_PLS
*.opin pulse
*.iopin VDD
*.iopin VSS
A1 net1 clk NULL ~RST_PLS NULL NULL ddflop
A2 net2 clk2 NULL ~RST_PLS NULL NULL ddflop
A3 net3 clk4 NULL ~RST_PLS NULL NULL ddflop
A4 net4 clk8 NULL ~RST_PLS NULL NULL ddflop
A5 [delayed clk64] net7 d_lut_sky130_fd_sc_hd__xor2_1
A9 net5 clk16 NULL ~RST_PLS NULL NULL ddflop
A10 net6 clk32 NULL ~RST_PLS NULL NULL ddflop
A6 clk64 clk NULL ~RST_PLS NULL NULL ddflop
A7 net7 ~clk NULL ~RST_PLS NULL NULL ddflop

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_clk] [clk] todig_1v8
AA2D2 [a_pulse] [pulse] todig_1v8
AA2D3 [a_VDD] [VDD] todig_1v8
AA2D4 [a_VSS] [VSS] todig_1v8
AA2D5 [a_RST_PLS] [RST_PLS] todig_1v8

.ends

.GLOBAL GND

* sky130_fd_sc_hd__dfrbp_1 IQ
* sky130_fd_sc_hd__xor2_1 (A&!B) | (!A&B)
.model d_lut_sky130_fd_sc_hd__xor2_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0110")
* sky130_fd_sc_hd__dfrtp_1 IQ
* sky130_fd_sc_hd__dfrtn_1 IQ
.end
