magic
tech sky130A
magscale 1 2
timestamp 1667492310
<< error_p >>
rect -125 1072 -67 1078
rect 67 1072 125 1078
rect -125 1038 -113 1072
rect 67 1038 79 1072
rect -125 1032 -67 1038
rect 67 1032 125 1038
rect -221 -1038 -163 -1032
rect -29 -1038 29 -1032
rect 163 -1038 221 -1032
rect -221 -1072 -209 -1038
rect -29 -1072 -17 -1038
rect 163 -1072 175 -1038
rect -221 -1078 -163 -1072
rect -29 -1078 29 -1072
rect 163 -1078 221 -1072
<< nmos >>
rect -207 -1000 -177 1000
rect -111 -1000 -81 1000
rect -15 -1000 15 1000
rect 81 -1000 111 1000
rect 177 -1000 207 1000
<< ndiff >>
rect -269 988 -207 1000
rect -269 -988 -257 988
rect -223 -988 -207 988
rect -269 -1000 -207 -988
rect -177 988 -111 1000
rect -177 -988 -161 988
rect -127 -988 -111 988
rect -177 -1000 -111 -988
rect -81 988 -15 1000
rect -81 -988 -65 988
rect -31 -988 -15 988
rect -81 -1000 -15 -988
rect 15 988 81 1000
rect 15 -988 31 988
rect 65 -988 81 988
rect 15 -1000 81 -988
rect 111 988 177 1000
rect 111 -988 127 988
rect 161 -988 177 988
rect 111 -1000 177 -988
rect 207 988 269 1000
rect 207 -988 223 988
rect 257 -988 269 988
rect 207 -1000 269 -988
<< ndiffc >>
rect -257 -988 -223 988
rect -161 -988 -127 988
rect -65 -988 -31 988
rect 31 -988 65 988
rect 127 -988 161 988
rect 223 -988 257 988
<< poly >>
rect -129 1072 -63 1088
rect -129 1038 -113 1072
rect -79 1038 -63 1072
rect -207 1000 -177 1026
rect -129 1022 -63 1038
rect 63 1072 129 1088
rect 63 1038 79 1072
rect 113 1038 129 1072
rect -111 1000 -81 1022
rect -15 1000 15 1026
rect 63 1022 129 1038
rect 81 1000 111 1022
rect 177 1000 207 1026
rect -207 -1022 -177 -1000
rect -225 -1038 -159 -1022
rect -111 -1026 -81 -1000
rect -15 -1022 15 -1000
rect -225 -1072 -209 -1038
rect -175 -1072 -159 -1038
rect -225 -1088 -159 -1072
rect -33 -1038 33 -1022
rect 81 -1026 111 -1000
rect 177 -1022 207 -1000
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect -33 -1088 33 -1072
rect 159 -1038 225 -1022
rect 159 -1072 175 -1038
rect 209 -1072 225 -1038
rect 159 -1088 225 -1072
<< polycont >>
rect -113 1038 -79 1072
rect 79 1038 113 1072
rect -209 -1072 -175 -1038
rect -17 -1072 17 -1038
rect 175 -1072 209 -1038
<< locali >>
rect -129 1038 -113 1072
rect -79 1038 -63 1072
rect 63 1038 79 1072
rect 113 1038 129 1072
rect -257 988 -223 1004
rect -257 -1004 -223 -988
rect -161 988 -127 1004
rect -161 -1004 -127 -988
rect -65 988 -31 1004
rect -65 -1004 -31 -988
rect 31 988 65 1004
rect 31 -1004 65 -988
rect 127 988 161 1004
rect 127 -1004 161 -988
rect 223 988 257 1004
rect 223 -1004 257 -988
rect -225 -1072 -209 -1038
rect -175 -1072 -159 -1038
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect 159 -1072 175 -1038
rect 209 -1072 225 -1038
<< viali >>
rect -113 1038 -79 1072
rect 79 1038 113 1072
rect -257 -971 -223 17
rect -161 -988 -127 988
rect -65 -971 -31 17
rect 31 -988 65 988
rect 127 -971 161 17
rect 223 -988 257 988
rect -209 -1072 -175 -1038
rect -17 -1072 17 -1038
rect 175 -1072 209 -1038
<< metal1 >>
rect -125 1072 -67 1078
rect -125 1038 -113 1072
rect -79 1038 -67 1072
rect -125 1032 -67 1038
rect 67 1072 125 1078
rect 67 1038 79 1072
rect 113 1038 125 1072
rect 67 1032 125 1038
rect -167 988 -121 1000
rect -263 17 -217 29
rect -263 -971 -257 17
rect -223 -971 -217 17
rect -263 -983 -217 -971
rect -167 -988 -161 988
rect -127 -988 -121 988
rect 25 988 71 1000
rect -71 17 -25 29
rect -71 -971 -65 17
rect -31 -971 -25 17
rect -71 -983 -25 -971
rect -167 -1000 -121 -988
rect 25 -988 31 988
rect 65 -988 71 988
rect 217 988 263 1000
rect 121 17 167 29
rect 121 -971 127 17
rect 161 -971 167 17
rect 121 -983 167 -971
rect 25 -1000 71 -988
rect 217 -988 223 988
rect 257 -988 263 988
rect 217 -1000 263 -988
rect -221 -1038 -163 -1032
rect -221 -1072 -209 -1038
rect -175 -1072 -163 -1038
rect -221 -1078 -163 -1072
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect 17 -1072 29 -1038
rect -29 -1078 29 -1072
rect 163 -1038 221 -1032
rect 163 -1072 175 -1038
rect 209 -1072 221 -1038
rect 163 -1078 221 -1072
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn +50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
