magic
tech sky130A
magscale 1 2
timestamp 1666302571
<< metal3 >>
rect -3928 17972 -3156 18000
rect -3928 13738 -3240 17972
rect -3176 13738 -3156 17972
rect -3928 13710 -3156 13738
rect -2916 17972 -2144 18000
rect -2916 13738 -2228 17972
rect -2164 13738 -2144 17972
rect -2916 13710 -2144 13738
rect -1904 17972 -1132 18000
rect -1904 13738 -1216 17972
rect -1152 13738 -1132 17972
rect -1904 13710 -1132 13738
rect -892 17972 -120 18000
rect -892 13738 -204 17972
rect -140 13738 -120 17972
rect -892 13710 -120 13738
rect 120 17972 892 18000
rect 120 13738 808 17972
rect 872 13738 892 17972
rect 120 13710 892 13738
rect 1132 17972 1904 18000
rect 1132 13738 1820 17972
rect 1884 13738 1904 17972
rect 1132 13710 1904 13738
rect 2144 17972 2916 18000
rect 2144 13738 2832 17972
rect 2896 13738 2916 17972
rect 2144 13710 2916 13738
rect 3156 17972 3928 18000
rect 3156 13738 3844 17972
rect 3908 13738 3928 17972
rect 3156 13710 3928 13738
rect -3928 13442 -3156 13470
rect -3928 9208 -3240 13442
rect -3176 9208 -3156 13442
rect -3928 9180 -3156 9208
rect -2916 13442 -2144 13470
rect -2916 9208 -2228 13442
rect -2164 9208 -2144 13442
rect -2916 9180 -2144 9208
rect -1904 13442 -1132 13470
rect -1904 9208 -1216 13442
rect -1152 9208 -1132 13442
rect -1904 9180 -1132 9208
rect -892 13442 -120 13470
rect -892 9208 -204 13442
rect -140 9208 -120 13442
rect -892 9180 -120 9208
rect 120 13442 892 13470
rect 120 9208 808 13442
rect 872 9208 892 13442
rect 120 9180 892 9208
rect 1132 13442 1904 13470
rect 1132 9208 1820 13442
rect 1884 9208 1904 13442
rect 1132 9180 1904 9208
rect 2144 13442 2916 13470
rect 2144 9208 2832 13442
rect 2896 9208 2916 13442
rect 2144 9180 2916 9208
rect 3156 13442 3928 13470
rect 3156 9208 3844 13442
rect 3908 9208 3928 13442
rect 3156 9180 3928 9208
rect -3928 8912 -3156 8940
rect -3928 4678 -3240 8912
rect -3176 4678 -3156 8912
rect -3928 4650 -3156 4678
rect -2916 8912 -2144 8940
rect -2916 4678 -2228 8912
rect -2164 4678 -2144 8912
rect -2916 4650 -2144 4678
rect -1904 8912 -1132 8940
rect -1904 4678 -1216 8912
rect -1152 4678 -1132 8912
rect -1904 4650 -1132 4678
rect -892 8912 -120 8940
rect -892 4678 -204 8912
rect -140 4678 -120 8912
rect -892 4650 -120 4678
rect 120 8912 892 8940
rect 120 4678 808 8912
rect 872 4678 892 8912
rect 120 4650 892 4678
rect 1132 8912 1904 8940
rect 1132 4678 1820 8912
rect 1884 4678 1904 8912
rect 1132 4650 1904 4678
rect 2144 8912 2916 8940
rect 2144 4678 2832 8912
rect 2896 4678 2916 8912
rect 2144 4650 2916 4678
rect 3156 8912 3928 8940
rect 3156 4678 3844 8912
rect 3908 4678 3928 8912
rect 3156 4650 3928 4678
rect -3928 4382 -3156 4410
rect -3928 148 -3240 4382
rect -3176 148 -3156 4382
rect -3928 120 -3156 148
rect -2916 4382 -2144 4410
rect -2916 148 -2228 4382
rect -2164 148 -2144 4382
rect -2916 120 -2144 148
rect -1904 4382 -1132 4410
rect -1904 148 -1216 4382
rect -1152 148 -1132 4382
rect -1904 120 -1132 148
rect -892 4382 -120 4410
rect -892 148 -204 4382
rect -140 148 -120 4382
rect -892 120 -120 148
rect 120 4382 892 4410
rect 120 148 808 4382
rect 872 148 892 4382
rect 120 120 892 148
rect 1132 4382 1904 4410
rect 1132 148 1820 4382
rect 1884 148 1904 4382
rect 1132 120 1904 148
rect 2144 4382 2916 4410
rect 2144 148 2832 4382
rect 2896 148 2916 4382
rect 2144 120 2916 148
rect 3156 4382 3928 4410
rect 3156 148 3844 4382
rect 3908 148 3928 4382
rect 3156 120 3928 148
rect -3928 -148 -3156 -120
rect -3928 -4382 -3240 -148
rect -3176 -4382 -3156 -148
rect -3928 -4410 -3156 -4382
rect -2916 -148 -2144 -120
rect -2916 -4382 -2228 -148
rect -2164 -4382 -2144 -148
rect -2916 -4410 -2144 -4382
rect -1904 -148 -1132 -120
rect -1904 -4382 -1216 -148
rect -1152 -4382 -1132 -148
rect -1904 -4410 -1132 -4382
rect -892 -148 -120 -120
rect -892 -4382 -204 -148
rect -140 -4382 -120 -148
rect -892 -4410 -120 -4382
rect 120 -148 892 -120
rect 120 -4382 808 -148
rect 872 -4382 892 -148
rect 120 -4410 892 -4382
rect 1132 -148 1904 -120
rect 1132 -4382 1820 -148
rect 1884 -4382 1904 -148
rect 1132 -4410 1904 -4382
rect 2144 -148 2916 -120
rect 2144 -4382 2832 -148
rect 2896 -4382 2916 -148
rect 2144 -4410 2916 -4382
rect 3156 -148 3928 -120
rect 3156 -4382 3844 -148
rect 3908 -4382 3928 -148
rect 3156 -4410 3928 -4382
rect -3928 -4678 -3156 -4650
rect -3928 -8912 -3240 -4678
rect -3176 -8912 -3156 -4678
rect -3928 -8940 -3156 -8912
rect -2916 -4678 -2144 -4650
rect -2916 -8912 -2228 -4678
rect -2164 -8912 -2144 -4678
rect -2916 -8940 -2144 -8912
rect -1904 -4678 -1132 -4650
rect -1904 -8912 -1216 -4678
rect -1152 -8912 -1132 -4678
rect -1904 -8940 -1132 -8912
rect -892 -4678 -120 -4650
rect -892 -8912 -204 -4678
rect -140 -8912 -120 -4678
rect -892 -8940 -120 -8912
rect 120 -4678 892 -4650
rect 120 -8912 808 -4678
rect 872 -8912 892 -4678
rect 120 -8940 892 -8912
rect 1132 -4678 1904 -4650
rect 1132 -8912 1820 -4678
rect 1884 -8912 1904 -4678
rect 1132 -8940 1904 -8912
rect 2144 -4678 2916 -4650
rect 2144 -8912 2832 -4678
rect 2896 -8912 2916 -4678
rect 2144 -8940 2916 -8912
rect 3156 -4678 3928 -4650
rect 3156 -8912 3844 -4678
rect 3908 -8912 3928 -4678
rect 3156 -8940 3928 -8912
rect -3928 -9208 -3156 -9180
rect -3928 -13442 -3240 -9208
rect -3176 -13442 -3156 -9208
rect -3928 -13470 -3156 -13442
rect -2916 -9208 -2144 -9180
rect -2916 -13442 -2228 -9208
rect -2164 -13442 -2144 -9208
rect -2916 -13470 -2144 -13442
rect -1904 -9208 -1132 -9180
rect -1904 -13442 -1216 -9208
rect -1152 -13442 -1132 -9208
rect -1904 -13470 -1132 -13442
rect -892 -9208 -120 -9180
rect -892 -13442 -204 -9208
rect -140 -13442 -120 -9208
rect -892 -13470 -120 -13442
rect 120 -9208 892 -9180
rect 120 -13442 808 -9208
rect 872 -13442 892 -9208
rect 120 -13470 892 -13442
rect 1132 -9208 1904 -9180
rect 1132 -13442 1820 -9208
rect 1884 -13442 1904 -9208
rect 1132 -13470 1904 -13442
rect 2144 -9208 2916 -9180
rect 2144 -13442 2832 -9208
rect 2896 -13442 2916 -9208
rect 2144 -13470 2916 -13442
rect 3156 -9208 3928 -9180
rect 3156 -13442 3844 -9208
rect 3908 -13442 3928 -9208
rect 3156 -13470 3928 -13442
rect -3928 -13738 -3156 -13710
rect -3928 -17972 -3240 -13738
rect -3176 -17972 -3156 -13738
rect -3928 -18000 -3156 -17972
rect -2916 -13738 -2144 -13710
rect -2916 -17972 -2228 -13738
rect -2164 -17972 -2144 -13738
rect -2916 -18000 -2144 -17972
rect -1904 -13738 -1132 -13710
rect -1904 -17972 -1216 -13738
rect -1152 -17972 -1132 -13738
rect -1904 -18000 -1132 -17972
rect -892 -13738 -120 -13710
rect -892 -17972 -204 -13738
rect -140 -17972 -120 -13738
rect -892 -18000 -120 -17972
rect 120 -13738 892 -13710
rect 120 -17972 808 -13738
rect 872 -17972 892 -13738
rect 120 -18000 892 -17972
rect 1132 -13738 1904 -13710
rect 1132 -17972 1820 -13738
rect 1884 -17972 1904 -13738
rect 1132 -18000 1904 -17972
rect 2144 -13738 2916 -13710
rect 2144 -17972 2832 -13738
rect 2896 -17972 2916 -13738
rect 2144 -18000 2916 -17972
rect 3156 -13738 3928 -13710
rect 3156 -17972 3844 -13738
rect 3908 -17972 3928 -13738
rect 3156 -18000 3928 -17972
<< via3 >>
rect -3240 13738 -3176 17972
rect -2228 13738 -2164 17972
rect -1216 13738 -1152 17972
rect -204 13738 -140 17972
rect 808 13738 872 17972
rect 1820 13738 1884 17972
rect 2832 13738 2896 17972
rect 3844 13738 3908 17972
rect -3240 9208 -3176 13442
rect -2228 9208 -2164 13442
rect -1216 9208 -1152 13442
rect -204 9208 -140 13442
rect 808 9208 872 13442
rect 1820 9208 1884 13442
rect 2832 9208 2896 13442
rect 3844 9208 3908 13442
rect -3240 4678 -3176 8912
rect -2228 4678 -2164 8912
rect -1216 4678 -1152 8912
rect -204 4678 -140 8912
rect 808 4678 872 8912
rect 1820 4678 1884 8912
rect 2832 4678 2896 8912
rect 3844 4678 3908 8912
rect -3240 148 -3176 4382
rect -2228 148 -2164 4382
rect -1216 148 -1152 4382
rect -204 148 -140 4382
rect 808 148 872 4382
rect 1820 148 1884 4382
rect 2832 148 2896 4382
rect 3844 148 3908 4382
rect -3240 -4382 -3176 -148
rect -2228 -4382 -2164 -148
rect -1216 -4382 -1152 -148
rect -204 -4382 -140 -148
rect 808 -4382 872 -148
rect 1820 -4382 1884 -148
rect 2832 -4382 2896 -148
rect 3844 -4382 3908 -148
rect -3240 -8912 -3176 -4678
rect -2228 -8912 -2164 -4678
rect -1216 -8912 -1152 -4678
rect -204 -8912 -140 -4678
rect 808 -8912 872 -4678
rect 1820 -8912 1884 -4678
rect 2832 -8912 2896 -4678
rect 3844 -8912 3908 -4678
rect -3240 -13442 -3176 -9208
rect -2228 -13442 -2164 -9208
rect -1216 -13442 -1152 -9208
rect -204 -13442 -140 -9208
rect 808 -13442 872 -9208
rect 1820 -13442 1884 -9208
rect 2832 -13442 2896 -9208
rect 3844 -13442 3908 -9208
rect -3240 -17972 -3176 -13738
rect -2228 -17972 -2164 -13738
rect -1216 -17972 -1152 -13738
rect -204 -17972 -140 -13738
rect 808 -17972 872 -13738
rect 1820 -17972 1884 -13738
rect 2832 -17972 2896 -13738
rect 3844 -17972 3908 -13738
<< mimcap >>
rect -3888 17920 -3488 17960
rect -3888 13790 -3848 17920
rect -3528 13790 -3488 17920
rect -3888 13750 -3488 13790
rect -2876 17920 -2476 17960
rect -2876 13790 -2836 17920
rect -2516 13790 -2476 17920
rect -2876 13750 -2476 13790
rect -1864 17920 -1464 17960
rect -1864 13790 -1824 17920
rect -1504 13790 -1464 17920
rect -1864 13750 -1464 13790
rect -852 17920 -452 17960
rect -852 13790 -812 17920
rect -492 13790 -452 17920
rect -852 13750 -452 13790
rect 160 17920 560 17960
rect 160 13790 200 17920
rect 520 13790 560 17920
rect 160 13750 560 13790
rect 1172 17920 1572 17960
rect 1172 13790 1212 17920
rect 1532 13790 1572 17920
rect 1172 13750 1572 13790
rect 2184 17920 2584 17960
rect 2184 13790 2224 17920
rect 2544 13790 2584 17920
rect 2184 13750 2584 13790
rect 3196 17920 3596 17960
rect 3196 13790 3236 17920
rect 3556 13790 3596 17920
rect 3196 13750 3596 13790
rect -3888 13390 -3488 13430
rect -3888 9260 -3848 13390
rect -3528 9260 -3488 13390
rect -3888 9220 -3488 9260
rect -2876 13390 -2476 13430
rect -2876 9260 -2836 13390
rect -2516 9260 -2476 13390
rect -2876 9220 -2476 9260
rect -1864 13390 -1464 13430
rect -1864 9260 -1824 13390
rect -1504 9260 -1464 13390
rect -1864 9220 -1464 9260
rect -852 13390 -452 13430
rect -852 9260 -812 13390
rect -492 9260 -452 13390
rect -852 9220 -452 9260
rect 160 13390 560 13430
rect 160 9260 200 13390
rect 520 9260 560 13390
rect 160 9220 560 9260
rect 1172 13390 1572 13430
rect 1172 9260 1212 13390
rect 1532 9260 1572 13390
rect 1172 9220 1572 9260
rect 2184 13390 2584 13430
rect 2184 9260 2224 13390
rect 2544 9260 2584 13390
rect 2184 9220 2584 9260
rect 3196 13390 3596 13430
rect 3196 9260 3236 13390
rect 3556 9260 3596 13390
rect 3196 9220 3596 9260
rect -3888 8860 -3488 8900
rect -3888 4730 -3848 8860
rect -3528 4730 -3488 8860
rect -3888 4690 -3488 4730
rect -2876 8860 -2476 8900
rect -2876 4730 -2836 8860
rect -2516 4730 -2476 8860
rect -2876 4690 -2476 4730
rect -1864 8860 -1464 8900
rect -1864 4730 -1824 8860
rect -1504 4730 -1464 8860
rect -1864 4690 -1464 4730
rect -852 8860 -452 8900
rect -852 4730 -812 8860
rect -492 4730 -452 8860
rect -852 4690 -452 4730
rect 160 8860 560 8900
rect 160 4730 200 8860
rect 520 4730 560 8860
rect 160 4690 560 4730
rect 1172 8860 1572 8900
rect 1172 4730 1212 8860
rect 1532 4730 1572 8860
rect 1172 4690 1572 4730
rect 2184 8860 2584 8900
rect 2184 4730 2224 8860
rect 2544 4730 2584 8860
rect 2184 4690 2584 4730
rect 3196 8860 3596 8900
rect 3196 4730 3236 8860
rect 3556 4730 3596 8860
rect 3196 4690 3596 4730
rect -3888 4330 -3488 4370
rect -3888 200 -3848 4330
rect -3528 200 -3488 4330
rect -3888 160 -3488 200
rect -2876 4330 -2476 4370
rect -2876 200 -2836 4330
rect -2516 200 -2476 4330
rect -2876 160 -2476 200
rect -1864 4330 -1464 4370
rect -1864 200 -1824 4330
rect -1504 200 -1464 4330
rect -1864 160 -1464 200
rect -852 4330 -452 4370
rect -852 200 -812 4330
rect -492 200 -452 4330
rect -852 160 -452 200
rect 160 4330 560 4370
rect 160 200 200 4330
rect 520 200 560 4330
rect 160 160 560 200
rect 1172 4330 1572 4370
rect 1172 200 1212 4330
rect 1532 200 1572 4330
rect 1172 160 1572 200
rect 2184 4330 2584 4370
rect 2184 200 2224 4330
rect 2544 200 2584 4330
rect 2184 160 2584 200
rect 3196 4330 3596 4370
rect 3196 200 3236 4330
rect 3556 200 3596 4330
rect 3196 160 3596 200
rect -3888 -200 -3488 -160
rect -3888 -4330 -3848 -200
rect -3528 -4330 -3488 -200
rect -3888 -4370 -3488 -4330
rect -2876 -200 -2476 -160
rect -2876 -4330 -2836 -200
rect -2516 -4330 -2476 -200
rect -2876 -4370 -2476 -4330
rect -1864 -200 -1464 -160
rect -1864 -4330 -1824 -200
rect -1504 -4330 -1464 -200
rect -1864 -4370 -1464 -4330
rect -852 -200 -452 -160
rect -852 -4330 -812 -200
rect -492 -4330 -452 -200
rect -852 -4370 -452 -4330
rect 160 -200 560 -160
rect 160 -4330 200 -200
rect 520 -4330 560 -200
rect 160 -4370 560 -4330
rect 1172 -200 1572 -160
rect 1172 -4330 1212 -200
rect 1532 -4330 1572 -200
rect 1172 -4370 1572 -4330
rect 2184 -200 2584 -160
rect 2184 -4330 2224 -200
rect 2544 -4330 2584 -200
rect 2184 -4370 2584 -4330
rect 3196 -200 3596 -160
rect 3196 -4330 3236 -200
rect 3556 -4330 3596 -200
rect 3196 -4370 3596 -4330
rect -3888 -4730 -3488 -4690
rect -3888 -8860 -3848 -4730
rect -3528 -8860 -3488 -4730
rect -3888 -8900 -3488 -8860
rect -2876 -4730 -2476 -4690
rect -2876 -8860 -2836 -4730
rect -2516 -8860 -2476 -4730
rect -2876 -8900 -2476 -8860
rect -1864 -4730 -1464 -4690
rect -1864 -8860 -1824 -4730
rect -1504 -8860 -1464 -4730
rect -1864 -8900 -1464 -8860
rect -852 -4730 -452 -4690
rect -852 -8860 -812 -4730
rect -492 -8860 -452 -4730
rect -852 -8900 -452 -8860
rect 160 -4730 560 -4690
rect 160 -8860 200 -4730
rect 520 -8860 560 -4730
rect 160 -8900 560 -8860
rect 1172 -4730 1572 -4690
rect 1172 -8860 1212 -4730
rect 1532 -8860 1572 -4730
rect 1172 -8900 1572 -8860
rect 2184 -4730 2584 -4690
rect 2184 -8860 2224 -4730
rect 2544 -8860 2584 -4730
rect 2184 -8900 2584 -8860
rect 3196 -4730 3596 -4690
rect 3196 -8860 3236 -4730
rect 3556 -8860 3596 -4730
rect 3196 -8900 3596 -8860
rect -3888 -9260 -3488 -9220
rect -3888 -13390 -3848 -9260
rect -3528 -13390 -3488 -9260
rect -3888 -13430 -3488 -13390
rect -2876 -9260 -2476 -9220
rect -2876 -13390 -2836 -9260
rect -2516 -13390 -2476 -9260
rect -2876 -13430 -2476 -13390
rect -1864 -9260 -1464 -9220
rect -1864 -13390 -1824 -9260
rect -1504 -13390 -1464 -9260
rect -1864 -13430 -1464 -13390
rect -852 -9260 -452 -9220
rect -852 -13390 -812 -9260
rect -492 -13390 -452 -9260
rect -852 -13430 -452 -13390
rect 160 -9260 560 -9220
rect 160 -13390 200 -9260
rect 520 -13390 560 -9260
rect 160 -13430 560 -13390
rect 1172 -9260 1572 -9220
rect 1172 -13390 1212 -9260
rect 1532 -13390 1572 -9260
rect 1172 -13430 1572 -13390
rect 2184 -9260 2584 -9220
rect 2184 -13390 2224 -9260
rect 2544 -13390 2584 -9260
rect 2184 -13430 2584 -13390
rect 3196 -9260 3596 -9220
rect 3196 -13390 3236 -9260
rect 3556 -13390 3596 -9260
rect 3196 -13430 3596 -13390
rect -3888 -13790 -3488 -13750
rect -3888 -17920 -3848 -13790
rect -3528 -17920 -3488 -13790
rect -3888 -17960 -3488 -17920
rect -2876 -13790 -2476 -13750
rect -2876 -17920 -2836 -13790
rect -2516 -17920 -2476 -13790
rect -2876 -17960 -2476 -17920
rect -1864 -13790 -1464 -13750
rect -1864 -17920 -1824 -13790
rect -1504 -17920 -1464 -13790
rect -1864 -17960 -1464 -17920
rect -852 -13790 -452 -13750
rect -852 -17920 -812 -13790
rect -492 -17920 -452 -13790
rect -852 -17960 -452 -17920
rect 160 -13790 560 -13750
rect 160 -17920 200 -13790
rect 520 -17920 560 -13790
rect 160 -17960 560 -17920
rect 1172 -13790 1572 -13750
rect 1172 -17920 1212 -13790
rect 1532 -17920 1572 -13790
rect 1172 -17960 1572 -17920
rect 2184 -13790 2584 -13750
rect 2184 -17920 2224 -13790
rect 2544 -17920 2584 -13790
rect 2184 -17960 2584 -17920
rect 3196 -13790 3596 -13750
rect 3196 -17920 3236 -13790
rect 3556 -17920 3596 -13790
rect 3196 -17960 3596 -17920
<< mimcapcontact >>
rect -3848 13790 -3528 17920
rect -2836 13790 -2516 17920
rect -1824 13790 -1504 17920
rect -812 13790 -492 17920
rect 200 13790 520 17920
rect 1212 13790 1532 17920
rect 2224 13790 2544 17920
rect 3236 13790 3556 17920
rect -3848 9260 -3528 13390
rect -2836 9260 -2516 13390
rect -1824 9260 -1504 13390
rect -812 9260 -492 13390
rect 200 9260 520 13390
rect 1212 9260 1532 13390
rect 2224 9260 2544 13390
rect 3236 9260 3556 13390
rect -3848 4730 -3528 8860
rect -2836 4730 -2516 8860
rect -1824 4730 -1504 8860
rect -812 4730 -492 8860
rect 200 4730 520 8860
rect 1212 4730 1532 8860
rect 2224 4730 2544 8860
rect 3236 4730 3556 8860
rect -3848 200 -3528 4330
rect -2836 200 -2516 4330
rect -1824 200 -1504 4330
rect -812 200 -492 4330
rect 200 200 520 4330
rect 1212 200 1532 4330
rect 2224 200 2544 4330
rect 3236 200 3556 4330
rect -3848 -4330 -3528 -200
rect -2836 -4330 -2516 -200
rect -1824 -4330 -1504 -200
rect -812 -4330 -492 -200
rect 200 -4330 520 -200
rect 1212 -4330 1532 -200
rect 2224 -4330 2544 -200
rect 3236 -4330 3556 -200
rect -3848 -8860 -3528 -4730
rect -2836 -8860 -2516 -4730
rect -1824 -8860 -1504 -4730
rect -812 -8860 -492 -4730
rect 200 -8860 520 -4730
rect 1212 -8860 1532 -4730
rect 2224 -8860 2544 -4730
rect 3236 -8860 3556 -4730
rect -3848 -13390 -3528 -9260
rect -2836 -13390 -2516 -9260
rect -1824 -13390 -1504 -9260
rect -812 -13390 -492 -9260
rect 200 -13390 520 -9260
rect 1212 -13390 1532 -9260
rect 2224 -13390 2544 -9260
rect 3236 -13390 3556 -9260
rect -3848 -17920 -3528 -13790
rect -2836 -17920 -2516 -13790
rect -1824 -17920 -1504 -13790
rect -812 -17920 -492 -13790
rect 200 -17920 520 -13790
rect 1212 -17920 1532 -13790
rect 2224 -17920 2544 -13790
rect 3236 -17920 3556 -13790
<< metal4 >>
rect -3740 17921 -3636 18120
rect -3256 17972 -3160 17988
rect -3849 17920 -3527 17921
rect -3849 13790 -3848 17920
rect -3528 13790 -3527 17920
rect -3849 13789 -3527 13790
rect -3740 13391 -3636 13789
rect -3256 13738 -3240 17972
rect -3176 13738 -3160 17972
rect -2728 17921 -2624 18120
rect -2244 17972 -2148 17988
rect -2837 17920 -2515 17921
rect -2837 13790 -2836 17920
rect -2516 13790 -2515 17920
rect -2837 13789 -2515 13790
rect -3256 13722 -3160 13738
rect -3256 13442 -3160 13458
rect -3849 13390 -3527 13391
rect -3849 9260 -3848 13390
rect -3528 9260 -3527 13390
rect -3849 9259 -3527 9260
rect -3740 8861 -3636 9259
rect -3256 9208 -3240 13442
rect -3176 9208 -3160 13442
rect -2728 13391 -2624 13789
rect -2244 13738 -2228 17972
rect -2164 13738 -2148 17972
rect -1716 17921 -1612 18120
rect -1232 17972 -1136 17988
rect -1825 17920 -1503 17921
rect -1825 13790 -1824 17920
rect -1504 13790 -1503 17920
rect -1825 13789 -1503 13790
rect -2244 13722 -2148 13738
rect -2244 13442 -2148 13458
rect -2837 13390 -2515 13391
rect -2837 9260 -2836 13390
rect -2516 9260 -2515 13390
rect -2837 9259 -2515 9260
rect -3256 9192 -3160 9208
rect -3256 8912 -3160 8928
rect -3849 8860 -3527 8861
rect -3849 4730 -3848 8860
rect -3528 4730 -3527 8860
rect -3849 4729 -3527 4730
rect -3740 4331 -3636 4729
rect -3256 4678 -3240 8912
rect -3176 4678 -3160 8912
rect -2728 8861 -2624 9259
rect -2244 9208 -2228 13442
rect -2164 9208 -2148 13442
rect -1716 13391 -1612 13789
rect -1232 13738 -1216 17972
rect -1152 13738 -1136 17972
rect -704 17921 -600 18120
rect -220 17972 -124 17988
rect -813 17920 -491 17921
rect -813 13790 -812 17920
rect -492 13790 -491 17920
rect -813 13789 -491 13790
rect -1232 13722 -1136 13738
rect -1232 13442 -1136 13458
rect -1825 13390 -1503 13391
rect -1825 9260 -1824 13390
rect -1504 9260 -1503 13390
rect -1825 9259 -1503 9260
rect -2244 9192 -2148 9208
rect -2244 8912 -2148 8928
rect -2837 8860 -2515 8861
rect -2837 4730 -2836 8860
rect -2516 4730 -2515 8860
rect -2837 4729 -2515 4730
rect -3256 4662 -3160 4678
rect -3256 4382 -3160 4398
rect -3849 4330 -3527 4331
rect -3849 200 -3848 4330
rect -3528 200 -3527 4330
rect -3849 199 -3527 200
rect -3740 -199 -3636 199
rect -3256 148 -3240 4382
rect -3176 148 -3160 4382
rect -2728 4331 -2624 4729
rect -2244 4678 -2228 8912
rect -2164 4678 -2148 8912
rect -1716 8861 -1612 9259
rect -1232 9208 -1216 13442
rect -1152 9208 -1136 13442
rect -704 13391 -600 13789
rect -220 13738 -204 17972
rect -140 13738 -124 17972
rect 308 17921 412 18120
rect 792 17972 888 17988
rect 199 17920 521 17921
rect 199 13790 200 17920
rect 520 13790 521 17920
rect 199 13789 521 13790
rect -220 13722 -124 13738
rect -220 13442 -124 13458
rect -813 13390 -491 13391
rect -813 9260 -812 13390
rect -492 9260 -491 13390
rect -813 9259 -491 9260
rect -1232 9192 -1136 9208
rect -1232 8912 -1136 8928
rect -1825 8860 -1503 8861
rect -1825 4730 -1824 8860
rect -1504 4730 -1503 8860
rect -1825 4729 -1503 4730
rect -2244 4662 -2148 4678
rect -2244 4382 -2148 4398
rect -2837 4330 -2515 4331
rect -2837 200 -2836 4330
rect -2516 200 -2515 4330
rect -2837 199 -2515 200
rect -3256 132 -3160 148
rect -3256 -148 -3160 -132
rect -3849 -200 -3527 -199
rect -3849 -4330 -3848 -200
rect -3528 -4330 -3527 -200
rect -3849 -4331 -3527 -4330
rect -3740 -4729 -3636 -4331
rect -3256 -4382 -3240 -148
rect -3176 -4382 -3160 -148
rect -2728 -199 -2624 199
rect -2244 148 -2228 4382
rect -2164 148 -2148 4382
rect -1716 4331 -1612 4729
rect -1232 4678 -1216 8912
rect -1152 4678 -1136 8912
rect -704 8861 -600 9259
rect -220 9208 -204 13442
rect -140 9208 -124 13442
rect 308 13391 412 13789
rect 792 13738 808 17972
rect 872 13738 888 17972
rect 1320 17921 1424 18120
rect 1804 17972 1900 17988
rect 1211 17920 1533 17921
rect 1211 13790 1212 17920
rect 1532 13790 1533 17920
rect 1211 13789 1533 13790
rect 792 13722 888 13738
rect 792 13442 888 13458
rect 199 13390 521 13391
rect 199 9260 200 13390
rect 520 9260 521 13390
rect 199 9259 521 9260
rect -220 9192 -124 9208
rect -220 8912 -124 8928
rect -813 8860 -491 8861
rect -813 4730 -812 8860
rect -492 4730 -491 8860
rect -813 4729 -491 4730
rect -1232 4662 -1136 4678
rect -1232 4382 -1136 4398
rect -1825 4330 -1503 4331
rect -1825 200 -1824 4330
rect -1504 200 -1503 4330
rect -1825 199 -1503 200
rect -2244 132 -2148 148
rect -2244 -148 -2148 -132
rect -2837 -200 -2515 -199
rect -2837 -4330 -2836 -200
rect -2516 -4330 -2515 -200
rect -2837 -4331 -2515 -4330
rect -3256 -4398 -3160 -4382
rect -3256 -4678 -3160 -4662
rect -3849 -4730 -3527 -4729
rect -3849 -8860 -3848 -4730
rect -3528 -8860 -3527 -4730
rect -3849 -8861 -3527 -8860
rect -3740 -9259 -3636 -8861
rect -3256 -8912 -3240 -4678
rect -3176 -8912 -3160 -4678
rect -2728 -4729 -2624 -4331
rect -2244 -4382 -2228 -148
rect -2164 -4382 -2148 -148
rect -1716 -199 -1612 199
rect -1232 148 -1216 4382
rect -1152 148 -1136 4382
rect -704 4331 -600 4729
rect -220 4678 -204 8912
rect -140 4678 -124 8912
rect 308 8861 412 9259
rect 792 9208 808 13442
rect 872 9208 888 13442
rect 1320 13391 1424 13789
rect 1804 13738 1820 17972
rect 1884 13738 1900 17972
rect 2332 17921 2436 18120
rect 2816 17972 2912 17988
rect 2223 17920 2545 17921
rect 2223 13790 2224 17920
rect 2544 13790 2545 17920
rect 2223 13789 2545 13790
rect 1804 13722 1900 13738
rect 1804 13442 1900 13458
rect 1211 13390 1533 13391
rect 1211 9260 1212 13390
rect 1532 9260 1533 13390
rect 1211 9259 1533 9260
rect 792 9192 888 9208
rect 792 8912 888 8928
rect 199 8860 521 8861
rect 199 4730 200 8860
rect 520 4730 521 8860
rect 199 4729 521 4730
rect -220 4662 -124 4678
rect -220 4382 -124 4398
rect -813 4330 -491 4331
rect -813 200 -812 4330
rect -492 200 -491 4330
rect -813 199 -491 200
rect -1232 132 -1136 148
rect -1232 -148 -1136 -132
rect -1825 -200 -1503 -199
rect -1825 -4330 -1824 -200
rect -1504 -4330 -1503 -200
rect -1825 -4331 -1503 -4330
rect -2244 -4398 -2148 -4382
rect -2244 -4678 -2148 -4662
rect -2837 -4730 -2515 -4729
rect -2837 -8860 -2836 -4730
rect -2516 -8860 -2515 -4730
rect -2837 -8861 -2515 -8860
rect -3256 -8928 -3160 -8912
rect -3256 -9208 -3160 -9192
rect -3849 -9260 -3527 -9259
rect -3849 -13390 -3848 -9260
rect -3528 -13390 -3527 -9260
rect -3849 -13391 -3527 -13390
rect -3740 -13789 -3636 -13391
rect -3256 -13442 -3240 -9208
rect -3176 -13442 -3160 -9208
rect -2728 -9259 -2624 -8861
rect -2244 -8912 -2228 -4678
rect -2164 -8912 -2148 -4678
rect -1716 -4729 -1612 -4331
rect -1232 -4382 -1216 -148
rect -1152 -4382 -1136 -148
rect -704 -199 -600 199
rect -220 148 -204 4382
rect -140 148 -124 4382
rect 308 4331 412 4729
rect 792 4678 808 8912
rect 872 4678 888 8912
rect 1320 8861 1424 9259
rect 1804 9208 1820 13442
rect 1884 9208 1900 13442
rect 2332 13391 2436 13789
rect 2816 13738 2832 17972
rect 2896 13738 2912 17972
rect 3344 17921 3448 18120
rect 3828 17972 3924 17988
rect 3235 17920 3557 17921
rect 3235 13790 3236 17920
rect 3556 13790 3557 17920
rect 3235 13789 3557 13790
rect 2816 13722 2912 13738
rect 2816 13442 2912 13458
rect 2223 13390 2545 13391
rect 2223 9260 2224 13390
rect 2544 9260 2545 13390
rect 2223 9259 2545 9260
rect 1804 9192 1900 9208
rect 1804 8912 1900 8928
rect 1211 8860 1533 8861
rect 1211 4730 1212 8860
rect 1532 4730 1533 8860
rect 1211 4729 1533 4730
rect 792 4662 888 4678
rect 792 4382 888 4398
rect 199 4330 521 4331
rect 199 200 200 4330
rect 520 200 521 4330
rect 199 199 521 200
rect -220 132 -124 148
rect -220 -148 -124 -132
rect -813 -200 -491 -199
rect -813 -4330 -812 -200
rect -492 -4330 -491 -200
rect -813 -4331 -491 -4330
rect -1232 -4398 -1136 -4382
rect -1232 -4678 -1136 -4662
rect -1825 -4730 -1503 -4729
rect -1825 -8860 -1824 -4730
rect -1504 -8860 -1503 -4730
rect -1825 -8861 -1503 -8860
rect -2244 -8928 -2148 -8912
rect -2244 -9208 -2148 -9192
rect -2837 -9260 -2515 -9259
rect -2837 -13390 -2836 -9260
rect -2516 -13390 -2515 -9260
rect -2837 -13391 -2515 -13390
rect -3256 -13458 -3160 -13442
rect -3256 -13738 -3160 -13722
rect -3849 -13790 -3527 -13789
rect -3849 -17920 -3848 -13790
rect -3528 -17920 -3527 -13790
rect -3849 -17921 -3527 -17920
rect -3740 -18120 -3636 -17921
rect -3256 -17972 -3240 -13738
rect -3176 -17972 -3160 -13738
rect -2728 -13789 -2624 -13391
rect -2244 -13442 -2228 -9208
rect -2164 -13442 -2148 -9208
rect -1716 -9259 -1612 -8861
rect -1232 -8912 -1216 -4678
rect -1152 -8912 -1136 -4678
rect -704 -4729 -600 -4331
rect -220 -4382 -204 -148
rect -140 -4382 -124 -148
rect 308 -199 412 199
rect 792 148 808 4382
rect 872 148 888 4382
rect 1320 4331 1424 4729
rect 1804 4678 1820 8912
rect 1884 4678 1900 8912
rect 2332 8861 2436 9259
rect 2816 9208 2832 13442
rect 2896 9208 2912 13442
rect 3344 13391 3448 13789
rect 3828 13738 3844 17972
rect 3908 13738 3924 17972
rect 3828 13722 3924 13738
rect 3828 13442 3924 13458
rect 3235 13390 3557 13391
rect 3235 9260 3236 13390
rect 3556 9260 3557 13390
rect 3235 9259 3557 9260
rect 2816 9192 2912 9208
rect 2816 8912 2912 8928
rect 2223 8860 2545 8861
rect 2223 4730 2224 8860
rect 2544 4730 2545 8860
rect 2223 4729 2545 4730
rect 1804 4662 1900 4678
rect 1804 4382 1900 4398
rect 1211 4330 1533 4331
rect 1211 200 1212 4330
rect 1532 200 1533 4330
rect 1211 199 1533 200
rect 792 132 888 148
rect 792 -148 888 -132
rect 199 -200 521 -199
rect 199 -4330 200 -200
rect 520 -4330 521 -200
rect 199 -4331 521 -4330
rect -220 -4398 -124 -4382
rect -220 -4678 -124 -4662
rect -813 -4730 -491 -4729
rect -813 -8860 -812 -4730
rect -492 -8860 -491 -4730
rect -813 -8861 -491 -8860
rect -1232 -8928 -1136 -8912
rect -1232 -9208 -1136 -9192
rect -1825 -9260 -1503 -9259
rect -1825 -13390 -1824 -9260
rect -1504 -13390 -1503 -9260
rect -1825 -13391 -1503 -13390
rect -2244 -13458 -2148 -13442
rect -2244 -13738 -2148 -13722
rect -2837 -13790 -2515 -13789
rect -2837 -17920 -2836 -13790
rect -2516 -17920 -2515 -13790
rect -2837 -17921 -2515 -17920
rect -3256 -17988 -3160 -17972
rect -2728 -18120 -2624 -17921
rect -2244 -17972 -2228 -13738
rect -2164 -17972 -2148 -13738
rect -1716 -13789 -1612 -13391
rect -1232 -13442 -1216 -9208
rect -1152 -13442 -1136 -9208
rect -704 -9259 -600 -8861
rect -220 -8912 -204 -4678
rect -140 -8912 -124 -4678
rect 308 -4729 412 -4331
rect 792 -4382 808 -148
rect 872 -4382 888 -148
rect 1320 -199 1424 199
rect 1804 148 1820 4382
rect 1884 148 1900 4382
rect 2332 4331 2436 4729
rect 2816 4678 2832 8912
rect 2896 4678 2912 8912
rect 3344 8861 3448 9259
rect 3828 9208 3844 13442
rect 3908 9208 3924 13442
rect 3828 9192 3924 9208
rect 3828 8912 3924 8928
rect 3235 8860 3557 8861
rect 3235 4730 3236 8860
rect 3556 4730 3557 8860
rect 3235 4729 3557 4730
rect 2816 4662 2912 4678
rect 2816 4382 2912 4398
rect 2223 4330 2545 4331
rect 2223 200 2224 4330
rect 2544 200 2545 4330
rect 2223 199 2545 200
rect 1804 132 1900 148
rect 1804 -148 1900 -132
rect 1211 -200 1533 -199
rect 1211 -4330 1212 -200
rect 1532 -4330 1533 -200
rect 1211 -4331 1533 -4330
rect 792 -4398 888 -4382
rect 792 -4678 888 -4662
rect 199 -4730 521 -4729
rect 199 -8860 200 -4730
rect 520 -8860 521 -4730
rect 199 -8861 521 -8860
rect -220 -8928 -124 -8912
rect -220 -9208 -124 -9192
rect -813 -9260 -491 -9259
rect -813 -13390 -812 -9260
rect -492 -13390 -491 -9260
rect -813 -13391 -491 -13390
rect -1232 -13458 -1136 -13442
rect -1232 -13738 -1136 -13722
rect -1825 -13790 -1503 -13789
rect -1825 -17920 -1824 -13790
rect -1504 -17920 -1503 -13790
rect -1825 -17921 -1503 -17920
rect -2244 -17988 -2148 -17972
rect -1716 -18120 -1612 -17921
rect -1232 -17972 -1216 -13738
rect -1152 -17972 -1136 -13738
rect -704 -13789 -600 -13391
rect -220 -13442 -204 -9208
rect -140 -13442 -124 -9208
rect 308 -9259 412 -8861
rect 792 -8912 808 -4678
rect 872 -8912 888 -4678
rect 1320 -4729 1424 -4331
rect 1804 -4382 1820 -148
rect 1884 -4382 1900 -148
rect 2332 -199 2436 199
rect 2816 148 2832 4382
rect 2896 148 2912 4382
rect 3344 4331 3448 4729
rect 3828 4678 3844 8912
rect 3908 4678 3924 8912
rect 3828 4662 3924 4678
rect 3828 4382 3924 4398
rect 3235 4330 3557 4331
rect 3235 200 3236 4330
rect 3556 200 3557 4330
rect 3235 199 3557 200
rect 2816 132 2912 148
rect 2816 -148 2912 -132
rect 2223 -200 2545 -199
rect 2223 -4330 2224 -200
rect 2544 -4330 2545 -200
rect 2223 -4331 2545 -4330
rect 1804 -4398 1900 -4382
rect 1804 -4678 1900 -4662
rect 1211 -4730 1533 -4729
rect 1211 -8860 1212 -4730
rect 1532 -8860 1533 -4730
rect 1211 -8861 1533 -8860
rect 792 -8928 888 -8912
rect 792 -9208 888 -9192
rect 199 -9260 521 -9259
rect 199 -13390 200 -9260
rect 520 -13390 521 -9260
rect 199 -13391 521 -13390
rect -220 -13458 -124 -13442
rect -220 -13738 -124 -13722
rect -813 -13790 -491 -13789
rect -813 -17920 -812 -13790
rect -492 -17920 -491 -13790
rect -813 -17921 -491 -17920
rect -1232 -17988 -1136 -17972
rect -704 -18120 -600 -17921
rect -220 -17972 -204 -13738
rect -140 -17972 -124 -13738
rect 308 -13789 412 -13391
rect 792 -13442 808 -9208
rect 872 -13442 888 -9208
rect 1320 -9259 1424 -8861
rect 1804 -8912 1820 -4678
rect 1884 -8912 1900 -4678
rect 2332 -4729 2436 -4331
rect 2816 -4382 2832 -148
rect 2896 -4382 2912 -148
rect 3344 -199 3448 199
rect 3828 148 3844 4382
rect 3908 148 3924 4382
rect 3828 132 3924 148
rect 3828 -148 3924 -132
rect 3235 -200 3557 -199
rect 3235 -4330 3236 -200
rect 3556 -4330 3557 -200
rect 3235 -4331 3557 -4330
rect 2816 -4398 2912 -4382
rect 2816 -4678 2912 -4662
rect 2223 -4730 2545 -4729
rect 2223 -8860 2224 -4730
rect 2544 -8860 2545 -4730
rect 2223 -8861 2545 -8860
rect 1804 -8928 1900 -8912
rect 1804 -9208 1900 -9192
rect 1211 -9260 1533 -9259
rect 1211 -13390 1212 -9260
rect 1532 -13390 1533 -9260
rect 1211 -13391 1533 -13390
rect 792 -13458 888 -13442
rect 792 -13738 888 -13722
rect 199 -13790 521 -13789
rect 199 -17920 200 -13790
rect 520 -17920 521 -13790
rect 199 -17921 521 -17920
rect -220 -17988 -124 -17972
rect 308 -18120 412 -17921
rect 792 -17972 808 -13738
rect 872 -17972 888 -13738
rect 1320 -13789 1424 -13391
rect 1804 -13442 1820 -9208
rect 1884 -13442 1900 -9208
rect 2332 -9259 2436 -8861
rect 2816 -8912 2832 -4678
rect 2896 -8912 2912 -4678
rect 3344 -4729 3448 -4331
rect 3828 -4382 3844 -148
rect 3908 -4382 3924 -148
rect 3828 -4398 3924 -4382
rect 3828 -4678 3924 -4662
rect 3235 -4730 3557 -4729
rect 3235 -8860 3236 -4730
rect 3556 -8860 3557 -4730
rect 3235 -8861 3557 -8860
rect 2816 -8928 2912 -8912
rect 2816 -9208 2912 -9192
rect 2223 -9260 2545 -9259
rect 2223 -13390 2224 -9260
rect 2544 -13390 2545 -9260
rect 2223 -13391 2545 -13390
rect 1804 -13458 1900 -13442
rect 1804 -13738 1900 -13722
rect 1211 -13790 1533 -13789
rect 1211 -17920 1212 -13790
rect 1532 -17920 1533 -13790
rect 1211 -17921 1533 -17920
rect 792 -17988 888 -17972
rect 1320 -18120 1424 -17921
rect 1804 -17972 1820 -13738
rect 1884 -17972 1900 -13738
rect 2332 -13789 2436 -13391
rect 2816 -13442 2832 -9208
rect 2896 -13442 2912 -9208
rect 3344 -9259 3448 -8861
rect 3828 -8912 3844 -4678
rect 3908 -8912 3924 -4678
rect 3828 -8928 3924 -8912
rect 3828 -9208 3924 -9192
rect 3235 -9260 3557 -9259
rect 3235 -13390 3236 -9260
rect 3556 -13390 3557 -9260
rect 3235 -13391 3557 -13390
rect 2816 -13458 2912 -13442
rect 2816 -13738 2912 -13722
rect 2223 -13790 2545 -13789
rect 2223 -17920 2224 -13790
rect 2544 -17920 2545 -13790
rect 2223 -17921 2545 -17920
rect 1804 -17988 1900 -17972
rect 2332 -18120 2436 -17921
rect 2816 -17972 2832 -13738
rect 2896 -17972 2912 -13738
rect 3344 -13789 3448 -13391
rect 3828 -13442 3844 -9208
rect 3908 -13442 3924 -9208
rect 3828 -13458 3924 -13442
rect 3828 -13738 3924 -13722
rect 3235 -13790 3557 -13789
rect 3235 -17920 3236 -13790
rect 3556 -17920 3557 -13790
rect 3235 -17921 3557 -17920
rect 2816 -17988 2912 -17972
rect 3344 -18120 3448 -17921
rect 3828 -17972 3844 -13738
rect 3908 -17972 3924 -13738
rect 3828 -17988 3924 -17972
<< properties >>
string FIXED_BBOX 3156 13710 3636 18000
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 8 ny 8 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
<< end >>
