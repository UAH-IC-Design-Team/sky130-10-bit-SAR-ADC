magic
tech sky130A
magscale 1 2
timestamp 1666918349
<< error_p >>
rect -29 2195 29 2201
rect -29 2161 -17 2195
rect -29 2155 29 2161
rect -29 1745 29 1751
rect -29 1711 -17 1745
rect -29 1705 29 1711
rect -29 1637 29 1643
rect -29 1603 -17 1637
rect -29 1597 29 1603
rect -29 1187 29 1193
rect -29 1153 -17 1187
rect -29 1147 29 1153
rect -29 1079 29 1085
rect -29 1045 -17 1079
rect -29 1039 29 1045
rect -29 629 29 635
rect -29 595 -17 629
rect -29 589 29 595
rect -29 521 29 527
rect -29 487 -17 521
rect -29 481 29 487
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -487 29 -481
rect -29 -521 -17 -487
rect -29 -527 29 -521
rect -29 -595 29 -589
rect -29 -629 -17 -595
rect -29 -635 29 -629
rect -29 -1045 29 -1039
rect -29 -1079 -17 -1045
rect -29 -1085 29 -1079
rect -29 -1153 29 -1147
rect -29 -1187 -17 -1153
rect -29 -1193 29 -1187
rect -29 -1603 29 -1597
rect -29 -1637 -17 -1603
rect -29 -1643 29 -1637
rect -29 -1711 29 -1705
rect -29 -1745 -17 -1711
rect -29 -1751 29 -1745
rect -29 -2161 29 -2155
rect -29 -2195 -17 -2161
rect -29 -2201 29 -2195
<< nwell >>
rect -211 -2333 211 2333
<< pmos >>
rect -15 1792 15 2114
rect -15 1234 15 1556
rect -15 676 15 998
rect -15 118 15 440
rect -15 -440 15 -118
rect -15 -998 15 -676
rect -15 -1556 15 -1234
rect -15 -2114 15 -1792
<< pdiff >>
rect -73 2102 -15 2114
rect -73 1804 -61 2102
rect -27 1804 -15 2102
rect -73 1792 -15 1804
rect 15 2102 73 2114
rect 15 1804 27 2102
rect 61 1804 73 2102
rect 15 1792 73 1804
rect -73 1544 -15 1556
rect -73 1246 -61 1544
rect -27 1246 -15 1544
rect -73 1234 -15 1246
rect 15 1544 73 1556
rect 15 1246 27 1544
rect 61 1246 73 1544
rect 15 1234 73 1246
rect -73 986 -15 998
rect -73 688 -61 986
rect -27 688 -15 986
rect -73 676 -15 688
rect 15 986 73 998
rect 15 688 27 986
rect 61 688 73 986
rect 15 676 73 688
rect -73 428 -15 440
rect -73 130 -61 428
rect -27 130 -15 428
rect -73 118 -15 130
rect 15 428 73 440
rect 15 130 27 428
rect 61 130 73 428
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -428 -61 -130
rect -27 -428 -15 -130
rect -73 -440 -15 -428
rect 15 -130 73 -118
rect 15 -428 27 -130
rect 61 -428 73 -130
rect 15 -440 73 -428
rect -73 -688 -15 -676
rect -73 -986 -61 -688
rect -27 -986 -15 -688
rect -73 -998 -15 -986
rect 15 -688 73 -676
rect 15 -986 27 -688
rect 61 -986 73 -688
rect 15 -998 73 -986
rect -73 -1246 -15 -1234
rect -73 -1544 -61 -1246
rect -27 -1544 -15 -1246
rect -73 -1556 -15 -1544
rect 15 -1246 73 -1234
rect 15 -1544 27 -1246
rect 61 -1544 73 -1246
rect 15 -1556 73 -1544
rect -73 -1804 -15 -1792
rect -73 -2102 -61 -1804
rect -27 -2102 -15 -1804
rect -73 -2114 -15 -2102
rect 15 -1804 73 -1792
rect 15 -2102 27 -1804
rect 61 -2102 73 -1804
rect 15 -2114 73 -2102
<< pdiffc >>
rect -61 1804 -27 2102
rect 27 1804 61 2102
rect -61 1246 -27 1544
rect 27 1246 61 1544
rect -61 688 -27 986
rect 27 688 61 986
rect -61 130 -27 428
rect 27 130 61 428
rect -61 -428 -27 -130
rect 27 -428 61 -130
rect -61 -986 -27 -688
rect 27 -986 61 -688
rect -61 -1544 -27 -1246
rect 27 -1544 61 -1246
rect -61 -2102 -27 -1804
rect 27 -2102 61 -1804
<< nsubdiff >>
rect -175 2263 -79 2297
rect 79 2263 175 2297
rect -175 2201 -141 2263
rect 141 2201 175 2263
rect -175 -2263 -141 -2201
rect 141 -2263 175 -2201
rect -175 -2297 -79 -2263
rect 79 -2297 175 -2263
<< nsubdiffcont >>
rect -79 2263 79 2297
rect -175 -2201 -141 2201
rect 141 -2201 175 2201
rect -79 -2297 79 -2263
<< poly >>
rect -33 2195 33 2211
rect -33 2161 -17 2195
rect 17 2161 33 2195
rect -33 2145 33 2161
rect -15 2114 15 2145
rect -15 1761 15 1792
rect -33 1745 33 1761
rect -33 1711 -17 1745
rect 17 1711 33 1745
rect -33 1695 33 1711
rect -33 1637 33 1653
rect -33 1603 -17 1637
rect 17 1603 33 1637
rect -33 1587 33 1603
rect -15 1556 15 1587
rect -15 1203 15 1234
rect -33 1187 33 1203
rect -33 1153 -17 1187
rect 17 1153 33 1187
rect -33 1137 33 1153
rect -33 1079 33 1095
rect -33 1045 -17 1079
rect 17 1045 33 1079
rect -33 1029 33 1045
rect -15 998 15 1029
rect -15 645 15 676
rect -33 629 33 645
rect -33 595 -17 629
rect 17 595 33 629
rect -33 579 33 595
rect -33 521 33 537
rect -33 487 -17 521
rect 17 487 33 521
rect -33 471 33 487
rect -15 440 15 471
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -471 15 -440
rect -33 -487 33 -471
rect -33 -521 -17 -487
rect 17 -521 33 -487
rect -33 -537 33 -521
rect -33 -595 33 -579
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -33 -645 33 -629
rect -15 -676 15 -645
rect -15 -1029 15 -998
rect -33 -1045 33 -1029
rect -33 -1079 -17 -1045
rect 17 -1079 33 -1045
rect -33 -1095 33 -1079
rect -33 -1153 33 -1137
rect -33 -1187 -17 -1153
rect 17 -1187 33 -1153
rect -33 -1203 33 -1187
rect -15 -1234 15 -1203
rect -15 -1587 15 -1556
rect -33 -1603 33 -1587
rect -33 -1637 -17 -1603
rect 17 -1637 33 -1603
rect -33 -1653 33 -1637
rect -33 -1711 33 -1695
rect -33 -1745 -17 -1711
rect 17 -1745 33 -1711
rect -33 -1761 33 -1745
rect -15 -1792 15 -1761
rect -15 -2145 15 -2114
rect -33 -2161 33 -2145
rect -33 -2195 -17 -2161
rect 17 -2195 33 -2161
rect -33 -2211 33 -2195
<< polycont >>
rect -17 2161 17 2195
rect -17 1711 17 1745
rect -17 1603 17 1637
rect -17 1153 17 1187
rect -17 1045 17 1079
rect -17 595 17 629
rect -17 487 17 521
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -521 17 -487
rect -17 -629 17 -595
rect -17 -1079 17 -1045
rect -17 -1187 17 -1153
rect -17 -1637 17 -1603
rect -17 -1745 17 -1711
rect -17 -2195 17 -2161
<< locali >>
rect -175 2263 -79 2297
rect 79 2263 175 2297
rect -175 2201 -141 2263
rect 141 2201 175 2263
rect -33 2161 -17 2195
rect 17 2161 33 2195
rect -61 2102 -27 2118
rect -61 1788 -27 1804
rect 27 2102 61 2118
rect 27 1788 61 1804
rect -33 1711 -17 1745
rect 17 1711 33 1745
rect -33 1603 -17 1637
rect 17 1603 33 1637
rect -61 1544 -27 1560
rect -61 1230 -27 1246
rect 27 1544 61 1560
rect 27 1230 61 1246
rect -33 1153 -17 1187
rect 17 1153 33 1187
rect -33 1045 -17 1079
rect 17 1045 33 1079
rect -61 986 -27 1002
rect -61 672 -27 688
rect 27 986 61 1002
rect 27 672 61 688
rect -33 595 -17 629
rect 17 595 33 629
rect -33 487 -17 521
rect 17 487 33 521
rect -61 428 -27 444
rect -61 114 -27 130
rect 27 428 61 444
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -444 -27 -428
rect 27 -130 61 -114
rect 27 -444 61 -428
rect -33 -521 -17 -487
rect 17 -521 33 -487
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -61 -688 -27 -672
rect -61 -1002 -27 -986
rect 27 -688 61 -672
rect 27 -1002 61 -986
rect -33 -1079 -17 -1045
rect 17 -1079 33 -1045
rect -33 -1187 -17 -1153
rect 17 -1187 33 -1153
rect -61 -1246 -27 -1230
rect -61 -1560 -27 -1544
rect 27 -1246 61 -1230
rect 27 -1560 61 -1544
rect -33 -1637 -17 -1603
rect 17 -1637 33 -1603
rect -33 -1745 -17 -1711
rect 17 -1745 33 -1711
rect -61 -1804 -27 -1788
rect -61 -2118 -27 -2102
rect 27 -1804 61 -1788
rect 27 -2118 61 -2102
rect -33 -2195 -17 -2161
rect 17 -2195 33 -2161
rect -175 -2263 -141 -2201
rect 141 -2263 175 -2201
rect -175 -2297 -79 -2263
rect 79 -2297 175 -2263
<< viali >>
rect -17 2161 17 2195
rect -61 1804 -27 2102
rect 27 1804 61 2102
rect -17 1711 17 1745
rect -17 1603 17 1637
rect -61 1246 -27 1544
rect 27 1246 61 1544
rect -17 1153 17 1187
rect -17 1045 17 1079
rect -61 688 -27 986
rect 27 688 61 986
rect -17 595 17 629
rect -17 487 17 521
rect -61 130 -27 428
rect 27 130 61 428
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -428 -27 -130
rect 27 -428 61 -130
rect -17 -521 17 -487
rect -17 -629 17 -595
rect -61 -986 -27 -688
rect 27 -986 61 -688
rect -17 -1079 17 -1045
rect -17 -1187 17 -1153
rect -61 -1544 -27 -1246
rect 27 -1544 61 -1246
rect -17 -1637 17 -1603
rect -17 -1745 17 -1711
rect -61 -2102 -27 -1804
rect 27 -2102 61 -1804
rect -17 -2195 17 -2161
<< metal1 >>
rect -29 2195 29 2201
rect -29 2161 -17 2195
rect 17 2161 29 2195
rect -29 2155 29 2161
rect -67 2102 -21 2114
rect -67 1804 -61 2102
rect -27 1804 -21 2102
rect -67 1792 -21 1804
rect 21 2102 67 2114
rect 21 1804 27 2102
rect 61 1804 67 2102
rect 21 1792 67 1804
rect -29 1745 29 1751
rect -29 1711 -17 1745
rect 17 1711 29 1745
rect -29 1705 29 1711
rect -29 1637 29 1643
rect -29 1603 -17 1637
rect 17 1603 29 1637
rect -29 1597 29 1603
rect -67 1544 -21 1556
rect -67 1246 -61 1544
rect -27 1246 -21 1544
rect -67 1234 -21 1246
rect 21 1544 67 1556
rect 21 1246 27 1544
rect 61 1246 67 1544
rect 21 1234 67 1246
rect -29 1187 29 1193
rect -29 1153 -17 1187
rect 17 1153 29 1187
rect -29 1147 29 1153
rect -29 1079 29 1085
rect -29 1045 -17 1079
rect 17 1045 29 1079
rect -29 1039 29 1045
rect -67 986 -21 998
rect -67 688 -61 986
rect -27 688 -21 986
rect -67 676 -21 688
rect 21 986 67 998
rect 21 688 27 986
rect 61 688 67 986
rect 21 676 67 688
rect -29 629 29 635
rect -29 595 -17 629
rect 17 595 29 629
rect -29 589 29 595
rect -29 521 29 527
rect -29 487 -17 521
rect 17 487 29 521
rect -29 481 29 487
rect -67 428 -21 440
rect -67 130 -61 428
rect -27 130 -21 428
rect -67 118 -21 130
rect 21 428 67 440
rect 21 130 27 428
rect 61 130 67 428
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -428 -61 -130
rect -27 -428 -21 -130
rect -67 -440 -21 -428
rect 21 -130 67 -118
rect 21 -428 27 -130
rect 61 -428 67 -130
rect 21 -440 67 -428
rect -29 -487 29 -481
rect -29 -521 -17 -487
rect 17 -521 29 -487
rect -29 -527 29 -521
rect -29 -595 29 -589
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -635 29 -629
rect -67 -688 -21 -676
rect -67 -986 -61 -688
rect -27 -986 -21 -688
rect -67 -998 -21 -986
rect 21 -688 67 -676
rect 21 -986 27 -688
rect 61 -986 67 -688
rect 21 -998 67 -986
rect -29 -1045 29 -1039
rect -29 -1079 -17 -1045
rect 17 -1079 29 -1045
rect -29 -1085 29 -1079
rect -29 -1153 29 -1147
rect -29 -1187 -17 -1153
rect 17 -1187 29 -1153
rect -29 -1193 29 -1187
rect -67 -1246 -21 -1234
rect -67 -1544 -61 -1246
rect -27 -1544 -21 -1246
rect -67 -1556 -21 -1544
rect 21 -1246 67 -1234
rect 21 -1544 27 -1246
rect 61 -1544 67 -1246
rect 21 -1556 67 -1544
rect -29 -1603 29 -1597
rect -29 -1637 -17 -1603
rect 17 -1637 29 -1603
rect -29 -1643 29 -1637
rect -29 -1711 29 -1705
rect -29 -1745 -17 -1711
rect 17 -1745 29 -1711
rect -29 -1751 29 -1745
rect -67 -1804 -21 -1792
rect -67 -2102 -61 -1804
rect -27 -2102 -21 -1804
rect -67 -2114 -21 -2102
rect 21 -1804 67 -1792
rect 21 -2102 27 -1804
rect 61 -2102 67 -1804
rect 21 -2114 67 -2102
rect -29 -2161 29 -2155
rect -29 -2195 -17 -2161
rect 17 -2195 29 -2161
rect -29 -2201 29 -2195
<< properties >>
string FIXED_BBOX -158 -2280 158 2280
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
