magic
tech sky130A
magscale 1 2
timestamp 1666555894
<< checkpaint >>
rect 3929 -1349 7847 1771
rect 9419 -1637 13337 1483
rect 18109 1043 21328 1051
rect 18109 -2069 21918 1043
rect 18770 -2117 21918 -2069
<< error_s >>
rect 1036 10791 1071 10825
rect 1037 10772 1071 10791
rect 867 10723 925 10729
rect 867 10689 879 10723
rect 867 10683 925 10689
rect 298 2915 333 2949
rect 721 2932 755 2950
rect 299 2896 333 2915
rect 129 2847 187 2853
rect 129 2813 141 2847
rect 129 2807 187 2813
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 2896
rect 352 2862 387 2896
rect 352 583 386 2862
rect 498 2794 556 2800
rect 498 2760 510 2794
rect 498 2754 556 2760
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 685 530 755 2932
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1056 477 1071 10772
rect 1090 10738 1125 10772
rect 1090 477 1124 10738
rect 1236 10670 1294 10676
rect 1236 10636 1248 10670
rect 1236 10630 1294 10636
rect 4749 4560 4784 4594
rect 4750 4541 4784 4560
rect 4580 4492 4638 4498
rect 4580 4458 4592 4492
rect 4580 4452 4638 4458
rect 4580 4042 4638 4048
rect 4580 4008 4592 4042
rect 4580 4002 4638 4008
rect 4580 3934 4638 3940
rect 4580 3900 4592 3934
rect 4580 3894 4638 3900
rect 4580 3484 4638 3490
rect 4580 3450 4592 3484
rect 4580 3444 4638 3450
rect 4580 3376 4638 3382
rect 4580 3342 4592 3376
rect 4580 3336 4638 3342
rect 4580 2926 4638 2932
rect 4580 2892 4592 2926
rect 4580 2886 4638 2892
rect 4580 2818 4638 2824
rect 1406 2769 1440 2787
rect 4580 2784 4592 2818
rect 4580 2778 4638 2784
rect 1406 2733 1476 2769
rect 1423 2699 1494 2733
rect 1774 2699 1809 2733
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1423 424 1493 2699
rect 1775 2680 1809 2699
rect 1605 2631 1663 2637
rect 1605 2597 1617 2631
rect 1605 2591 1663 2597
rect 1605 2181 1663 2187
rect 1605 2147 1617 2181
rect 1605 2141 1663 2147
rect 1605 2073 1663 2079
rect 1605 2039 1617 2073
rect 1605 2033 1663 2039
rect 1605 1623 1663 1629
rect 1605 1589 1617 1623
rect 1605 1583 1663 1589
rect 1605 1515 1663 1521
rect 1605 1481 1617 1515
rect 1605 1475 1663 1481
rect 1605 1065 1663 1071
rect 1605 1031 1617 1065
rect 1605 1025 1663 1031
rect 1605 957 1663 963
rect 1605 923 1617 957
rect 1605 917 1663 923
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1794 371 1809 2680
rect 1828 2646 1863 2680
rect 2143 2649 2178 2667
rect 2143 2646 2214 2649
rect 1828 371 1862 2646
rect 2144 2613 2214 2646
rect 1974 2578 2032 2584
rect 2161 2579 2232 2613
rect 1974 2544 1986 2578
rect 1974 2538 2032 2544
rect 1974 2128 2032 2134
rect 1974 2094 1986 2128
rect 1974 2088 2032 2094
rect 1974 2020 2032 2026
rect 1974 1986 1986 2020
rect 1974 1980 2032 1986
rect 1974 1570 2032 1576
rect 1974 1536 1986 1570
rect 1974 1530 2032 1536
rect 1974 1462 2032 1468
rect 1974 1428 1986 1462
rect 1974 1422 2032 1428
rect 1974 1012 2032 1018
rect 1974 978 1986 1012
rect 1974 972 2032 978
rect 1974 904 2032 910
rect 1974 870 1986 904
rect 1974 864 2032 870
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2161 318 2231 2579
rect 2443 2511 2501 2517
rect 2635 2511 2693 2517
rect 2443 2477 2455 2511
rect 2635 2477 2647 2511
rect 2443 2471 2501 2477
rect 2635 2471 2693 2477
rect 4580 2368 4638 2374
rect 4580 2334 4592 2368
rect 4580 2328 4638 2334
rect 4580 2260 4638 2266
rect 4580 2226 4592 2260
rect 4580 2220 4638 2226
rect 2905 1942 2939 1996
rect 2347 401 2405 407
rect 2539 401 2597 407
rect 2731 401 2789 407
rect 2347 367 2359 401
rect 2539 367 2551 401
rect 2731 367 2743 401
rect 2347 361 2405 367
rect 2539 361 2597 367
rect 2731 361 2789 367
rect 2161 282 2214 318
rect 2924 265 2939 1942
rect 2958 1908 2993 1942
rect 3273 1908 3308 1942
rect 2958 265 2992 1908
rect 3274 1889 3308 1908
rect 3104 1840 3162 1846
rect 3104 1806 3116 1840
rect 3104 1800 3162 1806
rect 3104 1548 3162 1554
rect 3104 1514 3116 1548
rect 3104 1508 3162 1514
rect 3104 1440 3162 1446
rect 3104 1406 3116 1440
rect 3104 1400 3162 1406
rect 3104 1148 3162 1154
rect 3104 1114 3116 1148
rect 3104 1108 3162 1114
rect 3104 1040 3162 1046
rect 3104 1006 3116 1040
rect 3104 1000 3162 1006
rect 3104 748 3162 754
rect 3104 714 3116 748
rect 3104 708 3162 714
rect 3104 640 3162 646
rect 3104 606 3116 640
rect 3104 600 3162 606
rect 3104 348 3162 354
rect 3104 314 3116 348
rect 3104 308 3162 314
rect 2958 231 2973 265
rect 3293 212 3308 1889
rect 3327 1855 3362 1889
rect 3642 1855 3677 1889
rect 3327 212 3361 1855
rect 3643 1836 3677 1855
rect 3473 1787 3531 1793
rect 3473 1753 3485 1787
rect 3473 1747 3531 1753
rect 3473 1495 3531 1501
rect 3473 1461 3485 1495
rect 3473 1455 3531 1461
rect 3473 1387 3531 1393
rect 3473 1353 3485 1387
rect 3473 1347 3531 1353
rect 3473 1095 3531 1101
rect 3473 1061 3485 1095
rect 3473 1055 3531 1061
rect 3473 987 3531 993
rect 3473 953 3485 987
rect 3473 947 3531 953
rect 3473 695 3531 701
rect 3473 661 3485 695
rect 3473 655 3531 661
rect 3473 587 3531 593
rect 3473 553 3485 587
rect 3473 547 3531 553
rect 3473 295 3531 301
rect 3473 261 3485 295
rect 3473 255 3531 261
rect 3327 178 3342 212
rect 3662 159 3677 1836
rect 3696 1802 3731 1836
rect 4011 1802 4046 1836
rect 4434 1819 4468 1837
rect 3696 159 3730 1802
rect 4012 1783 4046 1802
rect 3842 1734 3900 1740
rect 3842 1700 3854 1734
rect 3842 1694 3900 1700
rect 3842 1442 3900 1448
rect 3842 1408 3854 1442
rect 3842 1402 3900 1408
rect 3842 1334 3900 1340
rect 3842 1300 3854 1334
rect 3842 1294 3900 1300
rect 3842 1042 3900 1048
rect 3842 1008 3854 1042
rect 3842 1002 3900 1008
rect 3842 934 3900 940
rect 3842 900 3854 934
rect 3842 894 3900 900
rect 3842 642 3900 648
rect 3842 608 3854 642
rect 3842 602 3900 608
rect 3842 534 3900 540
rect 3842 500 3854 534
rect 3842 494 3900 500
rect 3842 242 3900 248
rect 3842 208 3854 242
rect 3842 202 3900 208
rect 3696 125 3711 159
rect 4031 106 4046 1783
rect 4065 1749 4100 1783
rect 4065 106 4099 1749
rect 4211 1681 4269 1687
rect 4211 1647 4223 1681
rect 4211 1641 4269 1647
rect 4211 1389 4269 1395
rect 4211 1355 4223 1389
rect 4211 1349 4269 1355
rect 4211 1281 4269 1287
rect 4211 1247 4223 1281
rect 4211 1241 4269 1247
rect 4211 989 4269 995
rect 4211 955 4223 989
rect 4211 949 4269 955
rect 4211 881 4269 887
rect 4211 847 4223 881
rect 4211 841 4269 847
rect 4211 589 4269 595
rect 4211 555 4223 589
rect 4211 549 4269 555
rect 4211 481 4269 487
rect 4211 447 4223 481
rect 4211 441 4269 447
rect 4211 189 4269 195
rect 4211 155 4223 189
rect 4211 149 4269 155
rect 4065 72 4080 106
rect 4398 53 4468 1819
rect 4580 1810 4638 1816
rect 4580 1776 4592 1810
rect 4580 1770 4638 1776
rect 4580 1702 4638 1708
rect 4580 1668 4592 1702
rect 4580 1662 4638 1668
rect 4580 1252 4638 1258
rect 4580 1218 4592 1252
rect 4580 1212 4638 1218
rect 4580 1144 4638 1150
rect 4580 1110 4592 1144
rect 4580 1104 4638 1110
rect 4580 694 4638 700
rect 4580 660 4592 694
rect 4580 654 4638 660
rect 4580 586 4638 592
rect 4580 552 4592 586
rect 4580 546 4638 552
rect 4580 136 4638 142
rect 4580 102 4592 136
rect 4580 96 4638 102
rect 4398 17 4451 53
rect 4769 0 4784 4541
rect 4803 4507 4838 4541
rect 4803 0 4837 4507
rect 4949 4439 5007 4445
rect 4949 4405 4961 4439
rect 4949 4399 5007 4405
rect 4949 3989 5007 3995
rect 4949 3955 4961 3989
rect 4949 3949 5007 3955
rect 4949 3881 5007 3887
rect 4949 3847 4961 3881
rect 4949 3841 5007 3847
rect 4949 3431 5007 3437
rect 4949 3397 4961 3431
rect 4949 3391 5007 3397
rect 4949 3323 5007 3329
rect 4949 3289 4961 3323
rect 4949 3283 5007 3289
rect 4949 2873 5007 2879
rect 4949 2839 4961 2873
rect 4949 2833 5007 2839
rect 4949 2765 5007 2771
rect 4949 2731 4961 2765
rect 4949 2725 5007 2731
rect 4949 2315 5007 2321
rect 4949 2281 4961 2315
rect 4949 2275 5007 2281
rect 4949 2207 5007 2213
rect 4949 2173 4961 2207
rect 4949 2167 5007 2173
rect 4949 1757 5007 1763
rect 4949 1723 4961 1757
rect 4949 1717 5007 1723
rect 4949 1649 5007 1655
rect 4949 1615 4961 1649
rect 4949 1609 5007 1615
rect 4949 1199 5007 1205
rect 4949 1165 4961 1199
rect 4949 1159 5007 1165
rect 4949 1091 5007 1097
rect 4949 1057 4961 1091
rect 4949 1051 5007 1057
rect 4949 641 5007 647
rect 4949 607 4961 641
rect 4949 601 5007 607
rect 4949 533 5007 539
rect 4949 499 4961 533
rect 4949 493 5007 499
rect 6863 124 6904 130
rect 4949 83 5007 89
rect 4949 49 4961 83
rect 7453 76 7466 108
rect 4949 43 5007 49
rect 4803 -34 4818 0
rect 8909 -20 8950 -14
rect 9499 -68 9512 -36
rect 12353 -164 12394 -158
rect 13533 -260 13574 -228
rect 15395 -404 15434 -372
rect 15801 -452 15842 -420
rect 16391 -500 16404 -468
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC1
timestamp 0
transform 1 0 5539 0 1 211
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC2
timestamp 0
transform 1 0 6238 0 1 211
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC3
timestamp 0
transform 1 0 11029 0 1 -77
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC4
timestamp 0
transform 1 0 11728 0 1 -77
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_4ZXHHB  XC5
timestamp 0
transform 1 0 18021 0 1 -409
box -450 -400 449 400
use sky130_fd_pr__cap_mim_m3_1_4ZXHHB  XC6
timestamp 0
transform 1 0 18920 0 1 -409
box -450 -400 449 400
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  XC7
timestamp 0
transform 1 0 19719 0 1 -509
box -350 -300 349 300
use sky130_fd_pr__pfet_01v8_XGA8MR  XM1
timestamp 0
transform 1 0 158 0 1 1766
box -211 -1219 211 1219
use sky130_fd_pr__pfet_01v8_XGA8MR  XM2
timestamp 0
transform 1 0 527 0 1 1713
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_SWP72P  XM3
timestamp 0
transform 1 0 896 0 1 5651
box -211 -5210 211 5210
use sky130_fd_pr__nfet_01v8_SWP72P  XM4
timestamp 0
transform 1 0 1265 0 1 5598
box -211 -5210 211 5210
use sky130_fd_pr__pfet_01v8_NF5RYF  XM5
timestamp 0
transform 1 0 1634 0 1 1552
box -211 -1217 211 1217
use sky130_fd_pr__pfet_01v8_NF5RYF  XM6
timestamp 0
transform 1 0 2003 0 1 1499
box -211 -1217 211 1217
use sky130_fd_pr__pfet_01v8_NF5ZBF  XM7
timestamp 0
transform 1 0 4609 0 1 2297
box -211 -2333 211 2333
use sky130_fd_pr__pfet_01v8_NF5ZBF  XM8
timestamp 0
transform 1 0 4978 0 1 2244
box -211 -2333 211 2333
use sky130_fd_pr__nfet_01v8_VJES5F  XM9
timestamp 0
transform 1 0 2568 0 1 1439
box -407 -1210 407 1210
use sky130_fd_pr__nfet_01v8_YBY378  XM11
timestamp 0
transform 1 0 3133 0 1 1077
box -211 -901 211 901
use sky130_fd_pr__nfet_01v8_YBY378  XM12
timestamp 0
transform 1 0 3502 0 1 1024
box -211 -901 211 901
use sky130_fd_pr__nfet_01v8_YBY378  XM13
timestamp 0
transform 1 0 3871 0 1 971
box -211 -901 211 901
use sky130_fd_pr__nfet_01v8_YBY378  XM14
timestamp 0
transform 1 0 4240 0 1 918
box -211 -901 211 901
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6587 0 1 -89
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6901 0 1 -137
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 7491 0 1 -185
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x4
timestamp 1662439860
transform 1 0 8633 0 1 -233
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x5
timestamp 1662439860
transform 1 0 8947 0 1 -281
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x6
timestamp 1662439860
transform 1 0 9537 0 1 -329
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x7
timestamp 1662439860
transform 1 0 12077 0 1 -377
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 12391 0 1 -425
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 13165 0 1 -473
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s15_1  x10
timestamp 1662439860
transform 1 0 13571 0 1 -521
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  x11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 14345 0 1 -569
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  x12
timestamp 1662439860
transform 1 0 15433 0 1 -665
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  x13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 15119 0 1 -617
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  x14
timestamp 1662439860
transform 1 0 15839 0 1 -713
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  x15
timestamp 1662439860
transform 1 0 16429 0 1 -761
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  x16
timestamp 1662439860
transform 1 0 20068 0 1 -809
box -38 -48 590 592
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin_p
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Out_n
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Vin_n
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Out_p
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 ext_clk
port 6 nsew
<< end >>
