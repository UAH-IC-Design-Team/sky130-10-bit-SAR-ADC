magic
tech sky130A
magscale 1 2
timestamp 1666724365
<< error_p >>
rect -119 62 -73 74
rect 73 62 119 74
rect -119 15 -113 62
rect 73 15 79 62
rect -119 3 -73 15
rect 73 3 119 15
rect -23 -15 23 -3
rect -23 -62 -17 -15
rect -23 -74 23 -62
<< nmos >>
rect -63 -91 -33 91
rect 33 -91 63 91
<< ndiff >>
rect -125 79 -63 91
rect -125 -79 -113 79
rect -79 -79 -63 79
rect -125 -91 -63 -79
rect -33 79 33 91
rect -33 -79 -17 79
rect 17 -79 33 79
rect -33 -91 33 -79
rect 63 79 125 91
rect 63 -79 79 79
rect 113 -79 125 79
rect 63 -91 125 -79
<< ndiffc >>
rect -113 -79 -79 79
rect -17 -79 17 79
rect 79 -79 113 79
<< poly >>
rect -63 91 -33 121
rect 33 91 63 121
rect -63 -113 -33 -91
rect 33 -113 63 -91
rect -85 -129 95 -113
rect -85 -163 -65 -129
rect -31 -163 25 -129
rect 59 -163 95 -129
rect -85 -179 95 -163
<< polycont >>
rect -65 -163 -31 -129
rect 25 -163 59 -129
<< locali >>
rect -113 79 -79 95
rect -113 -95 -79 -79
rect -17 79 17 95
rect -17 -95 17 -79
rect 79 79 113 95
rect 79 -95 113 -79
rect -85 -163 -65 -129
rect -31 -163 25 -129
rect 59 -163 95 -129
<< viali >>
rect -113 15 -79 62
rect -17 -62 17 -15
rect 79 15 113 62
rect -65 -163 -31 -129
rect 25 -163 59 -129
<< metal1 >>
rect -119 62 -73 74
rect -119 15 -113 62
rect -79 15 -73 62
rect -119 3 -73 15
rect 73 62 119 74
rect 73 15 79 62
rect 113 15 119 62
rect 73 3 119 15
rect -23 -15 23 -3
rect -23 -62 -17 -15
rect 17 -62 23 -15
rect -23 -74 23 -62
rect -85 -129 95 -123
rect -85 -163 -65 -129
rect -31 -163 25 -129
rect 59 -163 95 -129
rect -85 -169 95 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.91 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
