magic
tech sky130A
magscale 1 2
timestamp 1666918452
<< error_p >>
rect -29 5743 29 5749
rect -29 5709 -17 5743
rect -29 5703 29 5709
rect -29 4587 29 4593
rect -29 4553 -17 4587
rect -29 4547 29 4553
rect -29 3431 29 3437
rect -29 3397 -17 3431
rect -29 3391 29 3397
rect -29 2275 29 2281
rect -29 2241 -17 2275
rect -29 2235 29 2241
rect -29 1119 29 1125
rect -29 1085 -17 1119
rect -29 1079 29 1085
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -1193 29 -1187
rect -29 -1227 -17 -1193
rect -29 -1233 29 -1227
rect -29 -2349 29 -2343
rect -29 -2383 -17 -2349
rect -29 -2389 29 -2383
rect -29 -3505 29 -3499
rect -29 -3539 -17 -3505
rect -29 -3545 29 -3539
rect -29 -4661 29 -4655
rect -29 -4695 -17 -4661
rect -29 -4701 29 -4695
<< nmos >>
rect -15 4671 15 5671
rect -15 3515 15 4515
rect -15 2359 15 3359
rect -15 1203 15 2203
rect -15 47 15 1047
rect -15 -1109 15 -109
rect -15 -2265 15 -1265
rect -15 -3421 15 -2421
rect -15 -4577 15 -3577
rect -15 -5733 15 -4733
<< ndiff >>
rect -73 5659 -15 5671
rect -73 4683 -61 5659
rect -27 4683 -15 5659
rect -73 4671 -15 4683
rect 15 5659 73 5671
rect 15 4683 27 5659
rect 61 4683 73 5659
rect 15 4671 73 4683
rect -73 4503 -15 4515
rect -73 3527 -61 4503
rect -27 3527 -15 4503
rect -73 3515 -15 3527
rect 15 4503 73 4515
rect 15 3527 27 4503
rect 61 3527 73 4503
rect 15 3515 73 3527
rect -73 3347 -15 3359
rect -73 2371 -61 3347
rect -27 2371 -15 3347
rect -73 2359 -15 2371
rect 15 3347 73 3359
rect 15 2371 27 3347
rect 61 2371 73 3347
rect 15 2359 73 2371
rect -73 2191 -15 2203
rect -73 1215 -61 2191
rect -27 1215 -15 2191
rect -73 1203 -15 1215
rect 15 2191 73 2203
rect 15 1215 27 2191
rect 61 1215 73 2191
rect 15 1203 73 1215
rect -73 1035 -15 1047
rect -73 59 -61 1035
rect -27 59 -15 1035
rect -73 47 -15 59
rect 15 1035 73 1047
rect 15 59 27 1035
rect 61 59 73 1035
rect 15 47 73 59
rect -73 -121 -15 -109
rect -73 -1097 -61 -121
rect -27 -1097 -15 -121
rect -73 -1109 -15 -1097
rect 15 -121 73 -109
rect 15 -1097 27 -121
rect 61 -1097 73 -121
rect 15 -1109 73 -1097
rect -73 -1277 -15 -1265
rect -73 -2253 -61 -1277
rect -27 -2253 -15 -1277
rect -73 -2265 -15 -2253
rect 15 -1277 73 -1265
rect 15 -2253 27 -1277
rect 61 -2253 73 -1277
rect 15 -2265 73 -2253
rect -73 -2433 -15 -2421
rect -73 -3409 -61 -2433
rect -27 -3409 -15 -2433
rect -73 -3421 -15 -3409
rect 15 -2433 73 -2421
rect 15 -3409 27 -2433
rect 61 -3409 73 -2433
rect 15 -3421 73 -3409
rect -73 -3589 -15 -3577
rect -73 -4565 -61 -3589
rect -27 -4565 -15 -3589
rect -73 -4577 -15 -4565
rect 15 -3589 73 -3577
rect 15 -4565 27 -3589
rect 61 -4565 73 -3589
rect 15 -4577 73 -4565
rect -73 -4745 -15 -4733
rect -73 -5721 -61 -4745
rect -27 -5721 -15 -4745
rect -73 -5733 -15 -5721
rect 15 -4745 73 -4733
rect 15 -5721 27 -4745
rect 61 -5721 73 -4745
rect 15 -5733 73 -5721
<< ndiffc >>
rect -61 4683 -27 5659
rect 27 4683 61 5659
rect -61 3527 -27 4503
rect 27 3527 61 4503
rect -61 2371 -27 3347
rect 27 2371 61 3347
rect -61 1215 -27 2191
rect 27 1215 61 2191
rect -61 59 -27 1035
rect 27 59 61 1035
rect -61 -1097 -27 -121
rect 27 -1097 61 -121
rect -61 -2253 -27 -1277
rect 27 -2253 61 -1277
rect -61 -3409 -27 -2433
rect 27 -3409 61 -2433
rect -61 -4565 -27 -3589
rect 27 -4565 61 -3589
rect -61 -5721 -27 -4745
rect 27 -5721 61 -4745
<< poly >>
rect -33 5743 33 5759
rect -33 5709 -17 5743
rect 17 5709 33 5743
rect -33 5693 33 5709
rect -15 5671 15 5693
rect -15 4645 15 4671
rect -33 4587 33 4603
rect -33 4553 -17 4587
rect 17 4553 33 4587
rect -33 4537 33 4553
rect -15 4515 15 4537
rect -15 3489 15 3515
rect -33 3431 33 3447
rect -33 3397 -17 3431
rect 17 3397 33 3431
rect -33 3381 33 3397
rect -15 3359 15 3381
rect -15 2333 15 2359
rect -33 2275 33 2291
rect -33 2241 -17 2275
rect 17 2241 33 2275
rect -33 2225 33 2241
rect -15 2203 15 2225
rect -15 1177 15 1203
rect -33 1119 33 1135
rect -33 1085 -17 1119
rect 17 1085 33 1119
rect -33 1069 33 1085
rect -15 1047 15 1069
rect -15 21 15 47
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -1135 15 -1109
rect -33 -1193 33 -1177
rect -33 -1227 -17 -1193
rect 17 -1227 33 -1193
rect -33 -1243 33 -1227
rect -15 -1265 15 -1243
rect -15 -2291 15 -2265
rect -33 -2349 33 -2333
rect -33 -2383 -17 -2349
rect 17 -2383 33 -2349
rect -33 -2399 33 -2383
rect -15 -2421 15 -2399
rect -15 -3447 15 -3421
rect -33 -3505 33 -3489
rect -33 -3539 -17 -3505
rect 17 -3539 33 -3505
rect -33 -3555 33 -3539
rect -15 -3577 15 -3555
rect -15 -4603 15 -4577
rect -33 -4661 33 -4645
rect -33 -4695 -17 -4661
rect 17 -4695 33 -4661
rect -33 -4711 33 -4695
rect -15 -4733 15 -4711
rect -15 -5759 15 -5733
<< polycont >>
rect -17 5709 17 5743
rect -17 4553 17 4587
rect -17 3397 17 3431
rect -17 2241 17 2275
rect -17 1085 17 1119
rect -17 -71 17 -37
rect -17 -1227 17 -1193
rect -17 -2383 17 -2349
rect -17 -3539 17 -3505
rect -17 -4695 17 -4661
<< locali >>
rect -33 5709 -17 5743
rect 17 5709 33 5743
rect -61 5659 -27 5675
rect -61 4667 -27 4683
rect 27 5659 61 5675
rect 27 4667 61 4683
rect -33 4553 -17 4587
rect 17 4553 33 4587
rect -61 4503 -27 4519
rect -61 3511 -27 3527
rect 27 4503 61 4519
rect 27 3511 61 3527
rect -33 3397 -17 3431
rect 17 3397 33 3431
rect -61 3347 -27 3363
rect -61 2355 -27 2371
rect 27 3347 61 3363
rect 27 2355 61 2371
rect -33 2241 -17 2275
rect 17 2241 33 2275
rect -61 2191 -27 2207
rect -61 1199 -27 1215
rect 27 2191 61 2207
rect 27 1199 61 1215
rect -33 1085 -17 1119
rect 17 1085 33 1119
rect -61 1035 -27 1051
rect -61 43 -27 59
rect 27 1035 61 1051
rect 27 43 61 59
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -1113 -27 -1097
rect 27 -121 61 -105
rect 27 -1113 61 -1097
rect -33 -1227 -17 -1193
rect 17 -1227 33 -1193
rect -61 -1277 -27 -1261
rect -61 -2269 -27 -2253
rect 27 -1277 61 -1261
rect 27 -2269 61 -2253
rect -33 -2383 -17 -2349
rect 17 -2383 33 -2349
rect -61 -2433 -27 -2417
rect -61 -3425 -27 -3409
rect 27 -2433 61 -2417
rect 27 -3425 61 -3409
rect -33 -3539 -17 -3505
rect 17 -3539 33 -3505
rect -61 -3589 -27 -3573
rect -61 -4581 -27 -4565
rect 27 -3589 61 -3573
rect 27 -4581 61 -4565
rect -33 -4695 -17 -4661
rect 17 -4695 33 -4661
rect -61 -4745 -27 -4729
rect -61 -5737 -27 -5721
rect 27 -4745 61 -4729
rect 27 -5737 61 -5721
<< viali >>
rect -17 5709 17 5743
rect -61 4683 -27 5659
rect 27 4683 61 5659
rect -17 4553 17 4587
rect -61 3527 -27 4503
rect 27 3527 61 4503
rect -17 3397 17 3431
rect -61 2371 -27 3347
rect 27 2371 61 3347
rect -17 2241 17 2275
rect -61 1215 -27 2191
rect 27 1215 61 2191
rect -17 1085 17 1119
rect -61 59 -27 1035
rect 27 59 61 1035
rect -17 -71 17 -37
rect -61 -1097 -27 -121
rect 27 -1097 61 -121
rect -17 -1227 17 -1193
rect -61 -2253 -27 -1277
rect 27 -2253 61 -1277
rect -17 -2383 17 -2349
rect -61 -3409 -27 -2433
rect 27 -3409 61 -2433
rect -17 -3539 17 -3505
rect -61 -4565 -27 -3589
rect 27 -4565 61 -3589
rect -17 -4695 17 -4661
rect -61 -5721 -27 -4745
rect 27 -5721 61 -4745
<< metal1 >>
rect -29 5743 29 5749
rect -29 5709 -17 5743
rect 17 5709 29 5743
rect -29 5703 29 5709
rect -67 5659 -21 5671
rect -67 4683 -61 5659
rect -27 4683 -21 5659
rect -67 4671 -21 4683
rect 21 5659 67 5671
rect 21 4683 27 5659
rect 61 4683 67 5659
rect 21 4671 67 4683
rect -29 4587 29 4593
rect -29 4553 -17 4587
rect 17 4553 29 4587
rect -29 4547 29 4553
rect -67 4503 -21 4515
rect -67 3527 -61 4503
rect -27 3527 -21 4503
rect -67 3515 -21 3527
rect 21 4503 67 4515
rect 21 3527 27 4503
rect 61 3527 67 4503
rect 21 3515 67 3527
rect -29 3431 29 3437
rect -29 3397 -17 3431
rect 17 3397 29 3431
rect -29 3391 29 3397
rect -67 3347 -21 3359
rect -67 2371 -61 3347
rect -27 2371 -21 3347
rect -67 2359 -21 2371
rect 21 3347 67 3359
rect 21 2371 27 3347
rect 61 2371 67 3347
rect 21 2359 67 2371
rect -29 2275 29 2281
rect -29 2241 -17 2275
rect 17 2241 29 2275
rect -29 2235 29 2241
rect -67 2191 -21 2203
rect -67 1215 -61 2191
rect -27 1215 -21 2191
rect -67 1203 -21 1215
rect 21 2191 67 2203
rect 21 1215 27 2191
rect 61 1215 67 2191
rect 21 1203 67 1215
rect -29 1119 29 1125
rect -29 1085 -17 1119
rect 17 1085 29 1119
rect -29 1079 29 1085
rect -67 1035 -21 1047
rect -67 59 -61 1035
rect -27 59 -21 1035
rect -67 47 -21 59
rect 21 1035 67 1047
rect 21 59 27 1035
rect 61 59 67 1035
rect 21 47 67 59
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -1097 -61 -121
rect -27 -1097 -21 -121
rect -67 -1109 -21 -1097
rect 21 -121 67 -109
rect 21 -1097 27 -121
rect 61 -1097 67 -121
rect 21 -1109 67 -1097
rect -29 -1193 29 -1187
rect -29 -1227 -17 -1193
rect 17 -1227 29 -1193
rect -29 -1233 29 -1227
rect -67 -1277 -21 -1265
rect -67 -2253 -61 -1277
rect -27 -2253 -21 -1277
rect -67 -2265 -21 -2253
rect 21 -1277 67 -1265
rect 21 -2253 27 -1277
rect 61 -2253 67 -1277
rect 21 -2265 67 -2253
rect -29 -2349 29 -2343
rect -29 -2383 -17 -2349
rect 17 -2383 29 -2349
rect -29 -2389 29 -2383
rect -67 -2433 -21 -2421
rect -67 -3409 -61 -2433
rect -27 -3409 -21 -2433
rect -67 -3421 -21 -3409
rect 21 -2433 67 -2421
rect 21 -3409 27 -2433
rect 61 -3409 67 -2433
rect 21 -3421 67 -3409
rect -29 -3505 29 -3499
rect -29 -3539 -17 -3505
rect 17 -3539 29 -3505
rect -29 -3545 29 -3539
rect -67 -3589 -21 -3577
rect -67 -4565 -61 -3589
rect -27 -4565 -21 -3589
rect -67 -4577 -21 -4565
rect 21 -3589 67 -3577
rect 21 -4565 27 -3589
rect 61 -4565 67 -3589
rect 21 -4577 67 -4565
rect -29 -4661 29 -4655
rect -29 -4695 -17 -4661
rect 17 -4695 29 -4661
rect -29 -4701 29 -4695
rect -67 -4745 -21 -4733
rect -67 -5721 -61 -4745
rect -27 -5721 -21 -4745
rect -67 -5733 -21 -5721
rect 21 -4745 67 -4733
rect 21 -5721 27 -4745
rect 61 -5721 67 -4745
rect 21 -5733 67 -5721
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 10 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
