magic
tech sky130A
magscale 1 2
timestamp 1666650150
<< error_p >>
rect -1230 1200 -1170 3400
rect -1150 1200 -1090 3400
rect 1089 1200 1149 3400
rect 1169 1200 1229 3400
rect -1230 -1100 -1170 1100
rect -1150 -1100 -1090 1100
rect 1089 -1100 1149 1100
rect 1169 -1100 1229 1100
rect -1230 -3400 -1170 -1200
rect -1150 -3400 -1090 -1200
rect 1089 -3400 1149 -1200
rect 1169 -3400 1229 -1200
<< metal3 >>
rect -3469 3372 -1170 3400
rect -3469 1228 -1254 3372
rect -1190 1228 -1170 3372
rect -3469 1200 -1170 1228
rect -1150 3372 1149 3400
rect -1150 1228 1065 3372
rect 1129 1228 1149 3372
rect -1150 1200 1149 1228
rect 1169 3372 3468 3400
rect 1169 1228 3384 3372
rect 3448 1228 3468 3372
rect 1169 1200 3468 1228
rect -3469 1072 -1170 1100
rect -3469 -1072 -1254 1072
rect -1190 -1072 -1170 1072
rect -3469 -1100 -1170 -1072
rect -1150 1072 1149 1100
rect -1150 -1072 1065 1072
rect 1129 -1072 1149 1072
rect -1150 -1100 1149 -1072
rect 1169 1072 3468 1100
rect 1169 -1072 3384 1072
rect 3448 -1072 3468 1072
rect 1169 -1100 3468 -1072
rect -3469 -1228 -1170 -1200
rect -3469 -3372 -1254 -1228
rect -1190 -3372 -1170 -1228
rect -3469 -3400 -1170 -3372
rect -1150 -1228 1149 -1200
rect -1150 -3372 1065 -1228
rect 1129 -3372 1149 -1228
rect -1150 -3400 1149 -3372
rect 1169 -1228 3468 -1200
rect 1169 -3372 3384 -1228
rect 3448 -3372 3468 -1228
rect 1169 -3400 3468 -3372
<< via3 >>
rect -1254 1228 -1190 3372
rect 1065 1228 1129 3372
rect 3384 1228 3448 3372
rect -1254 -1072 -1190 1072
rect 1065 -1072 1129 1072
rect 3384 -1072 3448 1072
rect -1254 -3372 -1190 -1228
rect 1065 -3372 1129 -1228
rect 3384 -3372 3448 -1228
<< mimcap >>
rect -3369 3260 -1369 3300
rect -3369 1340 -3329 3260
rect -1409 1340 -1369 3260
rect -3369 1300 -1369 1340
rect -1050 3260 950 3300
rect -1050 1340 -1010 3260
rect 910 1340 950 3260
rect -1050 1300 950 1340
rect 1269 3260 3269 3300
rect 1269 1340 1309 3260
rect 3229 1340 3269 3260
rect 1269 1300 3269 1340
rect -3369 960 -1369 1000
rect -3369 -960 -3329 960
rect -1409 -960 -1369 960
rect -3369 -1000 -1369 -960
rect -1050 960 950 1000
rect -1050 -960 -1010 960
rect 910 -960 950 960
rect -1050 -1000 950 -960
rect 1269 960 3269 1000
rect 1269 -960 1309 960
rect 3229 -960 3269 960
rect 1269 -1000 3269 -960
rect -3369 -1340 -1369 -1300
rect -3369 -3260 -3329 -1340
rect -1409 -3260 -1369 -1340
rect -3369 -3300 -1369 -3260
rect -1050 -1340 950 -1300
rect -1050 -3260 -1010 -1340
rect 910 -3260 950 -1340
rect -1050 -3300 950 -3260
rect 1269 -1340 3269 -1300
rect 1269 -3260 1309 -1340
rect 3229 -3260 3269 -1340
rect 1269 -3300 3269 -3260
<< mimcapcontact >>
rect -3329 1340 -1409 3260
rect -1010 1340 910 3260
rect 1309 1340 3229 3260
rect -3329 -960 -1409 960
rect -1010 -960 910 960
rect 1309 -960 3229 960
rect -3329 -3260 -1409 -1340
rect -1010 -3260 910 -1340
rect 1309 -3260 3229 -1340
<< metal4 >>
rect -2421 3261 -2317 3450
rect -1301 3388 -1197 3450
rect -1301 3372 -1174 3388
rect -3330 3260 -1408 3261
rect -3330 1340 -3329 3260
rect -1409 1340 -1408 3260
rect -3330 1339 -1408 1340
rect -2421 961 -2317 1339
rect -1301 1228 -1254 3372
rect -1190 1228 -1174 3372
rect -102 3261 2 3450
rect 1018 3388 1122 3450
rect 1018 3372 1145 3388
rect -1011 3260 911 3261
rect -1011 1340 -1010 3260
rect 910 1340 911 3260
rect -1011 1339 911 1340
rect -1301 1212 -1174 1228
rect -1301 1088 -1197 1212
rect -1301 1072 -1174 1088
rect -3330 960 -1408 961
rect -3330 -960 -3329 960
rect -1409 -960 -1408 960
rect -3330 -961 -1408 -960
rect -2421 -1339 -2317 -961
rect -1301 -1072 -1254 1072
rect -1190 -1072 -1174 1072
rect -102 961 2 1339
rect 1018 1228 1065 3372
rect 1129 1228 1145 3372
rect 2217 3261 2321 3450
rect 3337 3388 3441 3450
rect 3337 3372 3464 3388
rect 1308 3260 3230 3261
rect 1308 1340 1309 3260
rect 3229 1340 3230 3260
rect 1308 1339 3230 1340
rect 1018 1212 1145 1228
rect 1018 1088 1122 1212
rect 1018 1072 1145 1088
rect -1011 960 911 961
rect -1011 -960 -1010 960
rect 910 -960 911 960
rect -1011 -961 911 -960
rect -1301 -1088 -1174 -1072
rect -1301 -1212 -1197 -1088
rect -1301 -1228 -1174 -1212
rect -3330 -1340 -1408 -1339
rect -3330 -3260 -3329 -1340
rect -1409 -3260 -1408 -1340
rect -3330 -3261 -1408 -3260
rect -2421 -3450 -2317 -3261
rect -1301 -3372 -1254 -1228
rect -1190 -3372 -1174 -1228
rect -102 -1339 2 -961
rect 1018 -1072 1065 1072
rect 1129 -1072 1145 1072
rect 2217 961 2321 1339
rect 3337 1228 3384 3372
rect 3448 1228 3464 3372
rect 3337 1212 3464 1228
rect 3337 1088 3441 1212
rect 3337 1072 3464 1088
rect 1308 960 3230 961
rect 1308 -960 1309 960
rect 3229 -960 3230 960
rect 1308 -961 3230 -960
rect 1018 -1088 1145 -1072
rect 1018 -1212 1122 -1088
rect 1018 -1228 1145 -1212
rect -1011 -1340 911 -1339
rect -1011 -3260 -1010 -1340
rect 910 -3260 911 -1340
rect -1011 -3261 911 -3260
rect -1301 -3388 -1174 -3372
rect -1301 -3450 -1197 -3388
rect -102 -3450 2 -3261
rect 1018 -3372 1065 -1228
rect 1129 -3372 1145 -1228
rect 2217 -1339 2321 -961
rect 3337 -1072 3384 1072
rect 3448 -1072 3464 1072
rect 3337 -1088 3464 -1072
rect 3337 -1212 3441 -1088
rect 3337 -1228 3464 -1212
rect 1308 -1340 3230 -1339
rect 1308 -3260 1309 -1340
rect 3229 -3260 3230 -1340
rect 1308 -3261 3230 -3260
rect 1018 -3388 1145 -3372
rect 1018 -3450 1122 -3388
rect 2217 -3450 2321 -3261
rect 3337 -3372 3384 -1228
rect 3448 -3372 3464 -1228
rect 3337 -3388 3464 -3372
rect 3337 -3450 3441 -3388
<< properties >>
string FIXED_BBOX 1169 1200 3369 3400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10 l 10 val 207.6 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
