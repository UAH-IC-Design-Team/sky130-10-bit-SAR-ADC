magic
tech sky130A
magscale 1 2
timestamp 1668283997
<< nwell >>
rect -5723822 -6577470 -5723501 -6577466
rect -5729320 -6577840 -5728999 -6577580
rect -5723822 -6577726 -5723499 -6577470
rect -5723820 -6577730 -5723499 -6577726
<< viali >>
rect -5729090 -6567670 -5729050 -6567530
rect -5726090 -6567840 -5726050 -6567710
rect -5723590 -6567850 -5723550 -6567710
rect -5729090 -6577770 -5729050 -6577630
rect -5723590 -6577650 -5723550 -6577520
rect -5726090 -6578030 -5726050 -6577890
<< metal1 >>
rect -5726580 -6566100 -5710100 -6566040
rect -5727300 -6566200 -5710100 -6566140
rect -5727840 -6566300 -5710100 -6566240
rect -5728540 -6566400 -5710100 -6566340
rect -5729080 -6566500 -5710100 -6566440
rect -5729780 -6566600 -5710100 -6566540
rect -5730320 -6566700 -5710100 -6566640
rect -5731020 -6566800 -5710100 -6566740
rect -5731560 -6566900 -5710100 -6566840
rect -5732260 -6567000 -5710100 -6566940
rect -5732800 -6567100 -5710100 -6567040
rect -5729100 -6567200 -5710100 -6567140
rect -5726100 -6567300 -5710100 -6567240
rect -5729370 -6567510 -5729270 -6567340
rect -5729370 -6567690 -5729360 -6567510
rect -5729280 -6567690 -5729270 -6567510
rect -5728830 -6567510 -5728730 -6567340
rect -5723600 -6567400 -5710100 -6567340
rect -5717780 -6567500 -5710100 -6567440
rect -5729370 -6567700 -5729270 -6567690
rect -5728830 -6567690 -5728820 -6567510
rect -5728740 -6567690 -5728730 -6567510
rect -5728830 -6567700 -5728730 -6567690
rect -5726330 -6567770 -5726230 -6567500
rect -5725790 -6567680 -5725690 -6567500
rect -5723830 -6567680 -5723730 -6567510
rect -5726430 -6567780 -5726230 -6567770
rect -5726430 -6567900 -5726420 -6567780
rect -5726310 -6567900 -5726230 -6567780
rect -5725790 -6567860 -5725780 -6567680
rect -5725700 -6567860 -5725690 -6567680
rect -5725790 -6567870 -5725690 -6567860
rect -5723910 -6567690 -5723730 -6567680
rect -5723910 -6567870 -5723900 -6567690
rect -5723810 -6567870 -5723730 -6567690
rect -5723290 -6567690 -5723190 -6567520
rect -5714880 -6567600 -5710100 -6567540
rect -5723910 -6567880 -5723730 -6567870
rect -5723290 -6567870 -5723280 -6567690
rect -5723200 -6567870 -5723190 -6567690
rect -5712380 -6567700 -5710100 -6567640
rect -5710760 -6567800 -5710100 -6567740
rect -5723290 -6567880 -5723190 -6567870
rect -5726430 -6567910 -5726230 -6567900
rect -5706344 -6568380 -5706268 -6568310
rect -5709300 -6570140 -5706700 -6570100
rect -5709300 -6570460 -5709260 -6570140
rect -5708040 -6570460 -5706700 -6570140
rect -5709300 -6570500 -5706700 -6570460
rect -5707660 -6570540 -5706700 -6570500
rect -5839600 -6571100 -5839510 -6571090
rect -5839600 -6571330 -5839590 -6571100
rect -5839520 -6571180 -5839510 -6571100
rect -5839520 -6571240 -5833280 -6571180
rect -5839520 -6571330 -5839510 -6571240
rect -5839600 -6571340 -5839510 -6571330
rect -5842270 -6571910 -5841950 -6571540
rect -5842100 -6572040 -5831500 -6572020
rect -5842100 -6572420 -5831880 -6572040
rect -5831520 -6572420 -5831500 -6572040
rect -5842100 -6572440 -5831500 -6572420
rect -5842100 -6572820 -5831500 -6572800
rect -5842100 -6573200 -5831880 -6572820
rect -5831520 -6573200 -5831500 -6572820
rect -5842100 -6573220 -5831500 -6573200
rect -5842270 -6573710 -5841950 -6573340
rect -5708600 -6574220 -5707700 -6574200
rect -5708600 -6574560 -5708560 -6574220
rect -5707720 -6574560 -5707700 -6574220
rect -5708600 -6574700 -5707700 -6574560
rect -5708600 -6574900 -5706700 -6574700
rect -5706341 -6576840 -5706262 -6576780
rect -5704960 -6577030 -5704840 -6576940
rect -5723930 -6577500 -5723730 -6577490
rect -5729330 -6577610 -5729230 -6577600
rect -5729330 -6577790 -5729320 -6577610
rect -5729240 -6577790 -5729230 -6577610
rect -5728790 -6577610 -5728680 -6577600
rect -5729330 -6577920 -5729230 -6577790
rect -5728790 -6577790 -5728780 -6577610
rect -5728690 -6577790 -5728680 -6577610
rect -5723930 -6577670 -5723920 -6577500
rect -5723810 -6577670 -5723730 -6577500
rect -5723300 -6577500 -5723190 -6577490
rect -5723930 -6577680 -5723730 -6577670
rect -5728790 -6577930 -5728680 -6577790
rect -5726340 -6577860 -5726240 -6577700
rect -5726420 -6577870 -5726240 -6577860
rect -5726420 -6578050 -5726410 -6577870
rect -5726310 -6578050 -5726240 -6577870
rect -5725800 -6577870 -5725700 -6577700
rect -5723830 -6577860 -5723730 -6577680
rect -5723300 -6577670 -5723290 -6577500
rect -5723200 -6577670 -5723190 -6577500
rect -5710760 -6577660 -5710100 -6577600
rect -5723300 -6577860 -5723190 -6577670
rect -5712380 -6577760 -5710100 -6577700
rect -5714880 -6577860 -5710100 -6577800
rect -5726420 -6578060 -5726240 -6578050
rect -5725800 -6578050 -5725790 -6577870
rect -5725710 -6578050 -5725700 -6577870
rect -5717780 -6577960 -5710100 -6577900
rect -5725800 -6578060 -5725700 -6578050
rect -5723600 -6578060 -5710100 -6578000
rect -5726100 -6578160 -5710100 -6578100
rect -5729100 -6578260 -5710100 -6578200
rect -5732800 -6578360 -5710100 -6578300
rect -5732260 -6578460 -5710100 -6578400
rect -5731560 -6578560 -5710100 -6578500
rect -5731020 -6578660 -5710100 -6578600
rect -5730320 -6578760 -5710100 -6578700
rect -5729780 -6578860 -5710100 -6578800
rect -5729080 -6578960 -5710100 -6578900
rect -5728540 -6579060 -5710100 -6579000
rect -5727840 -6579160 -5710100 -6579100
rect -5727300 -6579260 -5710100 -6579200
<< via1 >>
rect -5729360 -6567690 -5729280 -6567510
rect -5728820 -6567690 -5728740 -6567510
rect -5726420 -6567900 -5726310 -6567780
rect -5725780 -6567860 -5725700 -6567680
rect -5723900 -6567870 -5723810 -6567690
rect -5723280 -6567870 -5723200 -6567690
rect -5709260 -6570460 -5708040 -6570140
rect -5839590 -6571330 -5839520 -6571100
rect -5831880 -6572420 -5831520 -6572040
rect -5831880 -6573200 -5831520 -6572820
rect -5708560 -6574560 -5707720 -6574220
rect -5729320 -6577790 -5729240 -6577610
rect -5728780 -6577790 -5728690 -6577610
rect -5723920 -6577670 -5723810 -6577500
rect -5726410 -6578050 -5726310 -6577870
rect -5723290 -6577670 -5723200 -6577500
rect -5725790 -6578050 -5725710 -6577870
<< metal2 >>
rect -5729370 -6567510 -5729270 -6567500
rect -5729370 -6567690 -5729360 -6567510
rect -5729280 -6567690 -5729270 -6567510
rect -5729370 -6567700 -5729270 -6567690
rect -5728830 -6567510 -5728730 -6567500
rect -5728830 -6567690 -5728820 -6567510
rect -5728740 -6567690 -5728730 -6567510
rect -5728830 -6567700 -5728730 -6567690
rect -5725790 -6567680 -5725690 -6567670
rect -5726430 -6567780 -5726230 -6567770
rect -5726430 -6567900 -5726420 -6567780
rect -5726310 -6567900 -5726230 -6567780
rect -5725790 -6567860 -5725780 -6567680
rect -5725700 -6567860 -5725690 -6567680
rect -5725790 -6567870 -5725690 -6567860
rect -5723910 -6567690 -5723800 -6567680
rect -5723910 -6567870 -5723900 -6567690
rect -5723810 -6567870 -5723800 -6567690
rect -5723910 -6567880 -5723800 -6567870
rect -5723290 -6567690 -5723190 -6567680
rect -5723290 -6567870 -5723280 -6567690
rect -5723200 -6567870 -5723190 -6567690
rect -5723290 -6567880 -5723190 -6567870
rect -5726430 -6567910 -5726230 -6567900
rect -5709300 -6570140 -5708000 -6570100
rect -5709300 -6570460 -5709260 -6570140
rect -5708040 -6570460 -5708000 -6570140
rect -5709300 -6570500 -5708000 -6570460
rect -5831900 -6572040 -5831500 -6572020
rect -5831900 -6572420 -5831880 -6572040
rect -5831520 -6572420 -5831500 -6572040
rect -5831900 -6572440 -5831500 -6572420
rect -5831900 -6572820 -5831500 -6572800
rect -5831900 -6573200 -5831880 -6572820
rect -5831520 -6573200 -5831500 -6572820
rect -5831900 -6573220 -5831500 -6573200
rect -5708600 -6574220 -5707700 -6574200
rect -5708600 -6574560 -5708560 -6574220
rect -5707720 -6574560 -5707700 -6574220
rect -5708600 -6574600 -5707700 -6574560
rect -5723930 -6577500 -5723800 -6577490
rect -5729330 -6577610 -5729230 -6577600
rect -5729330 -6577790 -5729320 -6577610
rect -5729240 -6577790 -5729230 -6577610
rect -5729330 -6577800 -5729230 -6577790
rect -5728790 -6577610 -5728680 -6577600
rect -5728790 -6577790 -5728780 -6577610
rect -5728690 -6577790 -5728680 -6577610
rect -5723930 -6577670 -5723920 -6577500
rect -5723810 -6577670 -5723800 -6577500
rect -5723930 -6577680 -5723800 -6577670
rect -5723300 -6577500 -5723190 -6577490
rect -5723300 -6577670 -5723290 -6577500
rect -5723200 -6577670 -5723190 -6577500
rect -5723300 -6577680 -5723190 -6577670
rect -5728790 -6577800 -5728680 -6577790
rect -5726420 -6577870 -5726300 -6577860
rect -5726420 -6578050 -5726410 -6577870
rect -5726310 -6578050 -5726300 -6577870
rect -5726420 -6578060 -5726300 -6578050
rect -5725800 -6577870 -5725700 -6577860
rect -5725800 -6578050 -5725790 -6577870
rect -5725710 -6578050 -5725700 -6577870
rect -5725800 -6578060 -5725700 -6578050
<< via2 >>
rect -5729360 -6567690 -5729280 -6567510
rect -5728820 -6567690 -5728740 -6567510
rect -5726420 -6567900 -5726310 -6567780
rect -5725780 -6567860 -5725700 -6567680
rect -5723900 -6567870 -5723810 -6567690
rect -5723280 -6567870 -5723200 -6567690
rect -5709260 -6570460 -5708040 -6570140
rect -5831880 -6572420 -5831520 -6572040
rect -5840290 -6572790 -5840170 -6572450
rect -5839750 -6572790 -5839650 -6572450
rect -5707950 -6572790 -5707830 -6572440
rect -5831880 -6573200 -5831520 -6572820
rect -5708560 -6574560 -5707720 -6574220
rect -5708800 -6575300 -5708420 -6575160
rect -5729320 -6577790 -5729240 -6577610
rect -5728780 -6577790 -5728690 -6577610
rect -5723920 -6577670 -5723810 -6577500
rect -5723290 -6577670 -5723200 -6577500
rect -5726410 -6578050 -5726310 -6577870
rect -5725790 -6578050 -5725710 -6577870
<< metal3 >>
rect -5729370 -6567510 -5729270 -6567500
rect -5729370 -6567690 -5729360 -6567510
rect -5729280 -6567690 -5729270 -6567510
rect -5729370 -6567700 -5729270 -6567690
rect -5728830 -6567510 -5728730 -6567500
rect -5728830 -6567690 -5728820 -6567510
rect -5728740 -6567690 -5728730 -6567510
rect -5728830 -6567700 -5728730 -6567690
rect -5726430 -6567780 -5726230 -6567770
rect -5726430 -6567900 -5726420 -6567780
rect -5726310 -6567900 -5726230 -6567780
rect -5723910 -6567690 -5723800 -6567680
rect -5723910 -6567870 -5723900 -6567690
rect -5723810 -6567870 -5723800 -6567690
rect -5723910 -6567880 -5723800 -6567870
rect -5726430 -6567910 -5726230 -6567900
rect -5709300 -6570140 -5708000 -6570100
rect -5709300 -6570460 -5709260 -6570140
rect -5708040 -6570460 -5708000 -6570140
rect -5709300 -6570500 -5708000 -6570460
rect -5831900 -6572040 -5831500 -6572020
rect -5831900 -6572420 -5831880 -6572040
rect -5831520 -6572420 -5831500 -6572040
rect -5831900 -6572440 -5831500 -6572420
rect -5840300 -6572450 -5840160 -6572440
rect -5840300 -6572790 -5840290 -6572450
rect -5840170 -6572790 -5840160 -6572450
rect -5840300 -6572800 -5840160 -6572790
rect -5839760 -6572450 -5833600 -6572440
rect -5839760 -6572790 -5839750 -6572450
rect -5839650 -6572790 -5833600 -6572450
rect -5839760 -6572800 -5833600 -6572790
rect -5831900 -6572820 -5831500 -6572800
rect -5831900 -6573200 -5831880 -6572820
rect -5831520 -6573200 -5831500 -6572820
rect -5831900 -6573220 -5831500 -6573200
rect -5708600 -6574220 -5707700 -6574200
rect -5708600 -6574560 -5708560 -6574220
rect -5707720 -6574560 -5707700 -6574220
rect -5708600 -6574600 -5707700 -6574560
rect -5709800 -6575160 -5708400 -6575140
rect -5709800 -6575300 -5708800 -6575160
rect -5708420 -6575300 -5708400 -6575160
rect -5709800 -6575320 -5708400 -6575300
rect -5723930 -6577500 -5723800 -6577490
rect -5729330 -6577610 -5729230 -6577600
rect -5729330 -6577790 -5729320 -6577610
rect -5729240 -6577790 -5729230 -6577610
rect -5723930 -6577670 -5723920 -6577500
rect -5723810 -6577670 -5723800 -6577500
rect -5723930 -6577680 -5723800 -6577670
rect -5729330 -6577800 -5729230 -6577790
rect -5726420 -6577870 -5726300 -6577860
rect -5726420 -6578050 -5726410 -6577870
rect -5726310 -6578050 -5726300 -6577870
rect -5726420 -6578060 -5726300 -6578050
<< via3 >>
rect -5729360 -6567690 -5729280 -6567510
rect -5726420 -6567900 -5726310 -6567780
rect -5723900 -6567870 -5723810 -6567690
rect -5709260 -6570460 -5708040 -6570140
rect -5831880 -6572420 -5831520 -6572040
rect -5840290 -6572790 -5840170 -6572450
rect -5707950 -6572790 -5707830 -6572440
rect -5831880 -6573200 -5831520 -6572820
rect -5708560 -6574560 -5707720 -6574220
rect -5729320 -6577790 -5729240 -6577610
rect -5723920 -6577670 -5723810 -6577500
rect -5726410 -6578050 -5726310 -6577870
<< metal4 >>
rect -5709300 -6570140 -5708000 -6570100
rect -5709300 -6570460 -5709260 -6570140
rect -5708040 -6570460 -5708000 -6570140
rect -5709300 -6570500 -5708000 -6570460
rect -5831900 -6571500 -5716380 -6571100
rect -5831900 -6572040 -5831500 -6571500
rect -5831900 -6572420 -5831880 -6572040
rect -5831520 -6572420 -5831500 -6572040
rect -5831900 -6572440 -5831500 -6572420
rect -5709400 -6572440 -5707820 -6572420
rect -5840300 -6572450 -5833980 -6572440
rect -5840300 -6572790 -5840290 -6572450
rect -5840170 -6572790 -5833980 -6572450
rect -5840300 -6572800 -5833980 -6572790
rect -5709400 -6572790 -5707950 -6572440
rect -5707830 -6572790 -5707820 -6572440
rect -5709400 -6572800 -5707820 -6572790
rect -5831900 -6572820 -5831500 -6572800
rect -5831900 -6573200 -5831880 -6572820
rect -5831520 -6573200 -5831500 -6572820
rect -5831900 -6573700 -5831500 -6573200
rect -5831900 -6574100 -5716380 -6573700
rect -5708600 -6574220 -5707700 -6574200
rect -5708600 -6574560 -5708560 -6574220
rect -5707720 -6574560 -5707700 -6574220
rect -5708600 -6574600 -5707700 -6574560
<< via4 >>
rect -5709260 -6570460 -5708040 -6570140
rect -5711360 -6571460 -5710140 -6571140
rect -5711360 -6574060 -5710140 -6573740
rect -5708560 -6574560 -5707740 -6574240
<< metal5 >>
rect -5709300 -6570140 -5708000 -6570100
rect -5709300 -6570460 -5709260 -6570140
rect -5708040 -6570460 -5708000 -6570140
rect -5709300 -6570500 -5708000 -6570460
rect -5709300 -6571100 -5708700 -6570500
rect -5711400 -6571140 -5708700 -6571100
rect -5711400 -6571460 -5711360 -6571140
rect -5710140 -6571460 -5708700 -6571140
rect -5711400 -6571500 -5708700 -6571460
rect -5711400 -6573740 -5709400 -6573700
rect -5711400 -6574060 -5711360 -6573740
rect -5710140 -6574060 -5709400 -6573740
rect -5711400 -6574100 -5709400 -6574060
rect -5709920 -6574200 -5709400 -6574100
rect -5709920 -6574240 -5707700 -6574200
rect -5709920 -6574560 -5708560 -6574240
rect -5707740 -6574560 -5707700 -6574240
rect -5709920 -6574600 -5707700 -6574560
use bootstrapped_sampling_switch  bootstrapped_sampling_switch_0
timestamp 1668208340
transform 0 1 -5837200 1 0 -6579400
box -3600 -5100 17150 2800
use comparator  comparator_0
timestamp 1668204572
transform 0 -1 -5700550 1 0 -6584490
box 6930 4070 16410 8800
use dac  dac_0
timestamp 1668278360
transform 1 0 -5798000 0 1 -6624400
box -36000 33000 88600 70300
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 0 -1 -5728738 -1 0 -6577608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_1
timestamp 1662439860
transform 0 -1 -5723238 -1 0 -6567688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_2
timestamp 1662439860
transform 0 -1 -5728778 -1 0 -6567508
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_6
timestamp 1662439860
transform 0 -1 -5725748 -1 0 -6577868
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_7
timestamp 1662439860
transform 0 -1 -5725738 -1 0 -6567668
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_38
timestamp 1662439860
transform 0 -1 -5723238 -1 0 -6577498
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 0 -1 -5723238 -1 0 -6577760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1662439860
transform 0 -1 -5728738 -1 0 -6577870
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1662439860
transform 0 -1 -5725748 -1 0 -6577700
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1662439860
transform 0 -1 -5725738 -1 0 -6567510
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1662439860
transform 0 -1 -5728778 -1 0 -6567340
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1662439860
transform 0 -1 -5723238 -1 0 -6567520
box -38 -48 130 592
<< labels >>
rlabel metal4 -5709400 -6572800 -5707980 -6572420 1 VDD
port 1 n
rlabel metal1 -5842270 -6571910 -5841950 -6571540 1 V_in_p
port 2 n
rlabel metal3 -5709800 -6575320 -5708800 -6575140 1 VSS
port 3 n
rlabel metal1 -5842270 -6573710 -5841950 -6573340 1 V_in_n
port 4 n
rlabel metal1 -5706344 -6568380 -5706268 -6568310 1 comp_out_p
port 5 n
rlabel metal1 -5726580 -6566100 -5710100 -6566040 1 sw_sample_unbuf
port 6 n
rlabel metal1 -5704960 -6577030 -5704840 -6576940 1 comparator_clk
port 7 n
rlabel metal1 -5710760 -6577660 -5710100 -6577600 1 sw_sp_n9
port 8 n
rlabel metal1 -5723600 -6578060 -5710100 -6578000 1 sw_sp_n8
port 9 n
rlabel metal1 -5726100 -6578160 -5710100 -6578100 1 sw_sp_n7
port 10 n
rlabel metal1 -5729100 -6578260 -5710100 -6578200 1 sw_sp_n6
port 11 n
rlabel metal1 -5731020 -6578660 -5710100 -6578600 1 sw_sp_n5
port 12 n
rlabel metal1 -5730320 -6578760 -5710100 -6578700 1 sw_sp_n4
port 13 n
rlabel metal1 -5729780 -6578860 -5710100 -6578800 1 sw_sp_n3
port 14 n
rlabel metal1 -5727840 -6579160 -5710100 -6579100 1 sw_sp_n2
port 15 n
rlabel metal1 -5727300 -6579260 -5710100 -6579200 1 sw_sp_n1
port 16 n
rlabel metal1 -5710760 -6567800 -5710100 -6567740 1 sw_sp_p9
port 17 n
rlabel metal1 -5723600 -6567400 -5710100 -6567340 1 sw_sp_p8
port 18 n
rlabel metal1 -5726100 -6567300 -5710100 -6567240 1 sw_sp_p7
port 19 n
rlabel metal1 -5729100 -6567200 -5710100 -6567140 1 sw_sp_p6
port 20 n
rlabel metal1 -5731020 -6566800 -5710100 -6566740 1 sw_sp_p5
port 21 n
rlabel metal1 -5730320 -6566700 -5710100 -6566640 1 sw_sp_p4
port 22 n
rlabel metal1 -5729780 -6566600 -5710100 -6566540 1 sw_sp_p3
port 23 n
rlabel metal1 -5727840 -6566300 -5710100 -6566240 1 sw_sp_p2
port 24 n
rlabel metal1 -5727300 -6566200 -5710100 -6566140 1 sw_sp_p1
port 25 n
rlabel metal1 -5712380 -6577760 -5710100 -6577700 1 sw_n8
port 26 n
rlabel metal1 -5714880 -6577860 -5710100 -6577800 1 sw_n7
port 27 n
rlabel metal1 -5717780 -6577960 -5710100 -6577900 1 sw_n6
port 28 n
rlabel metal1 -5732800 -6578360 -5710100 -6578300 1 sw_n5
port 29 n
rlabel metal1 -5732260 -6578460 -5710100 -6578400 1 sw_n4
port 30 n
rlabel metal1 -5731560 -6578560 -5710100 -6578500 1 sw_n3
port 31 n
rlabel metal1 -5729080 -6578960 -5710100 -6578900 1 sw_n2
port 32 n
rlabel metal1 -5728540 -6579060 -5710100 -6579000 1 sw_n1
port 33 n
rlabel metal1 -5712380 -6567700 -5710100 -6567640 1 sw_p8
port 34 n
rlabel metal1 -5714880 -6567600 -5710100 -6567540 1 sw_p7
port 35 n
rlabel metal1 -5717780 -6567500 -5710100 -6567440 1 sw_p6
port 36 n
rlabel metal1 -5732800 -6567100 -5710100 -6567040 1 sw_p5
port 37 n
rlabel metal1 -5732260 -6567000 -5710100 -6566940 1 sw_p4
port 38 n
rlabel metal1 -5731560 -6566900 -5710100 -6566840 1 sw_p3
port 39 n
rlabel metal1 -5729080 -6566500 -5710100 -6566440 1 sw_p2
port 40 n
rlabel metal1 -5728540 -6566400 -5710100 -6566340 1 sw_p1
port 41 n
rlabel metal1 -5706341 -6576840 -5706262 -6576780 1 comp_out_n
port 42 n
<< end >>
