magic
tech sky130A
magscale 1 2
timestamp 1665882771
<< error_s >>
rect 671 1030 717 1042
rect 671 996 677 1030
rect 671 984 717 996
<< nwell >>
rect -300 910 730 1230
rect -300 900 240 910
<< psubdiff >>
rect 70 750 130 774
rect 70 626 130 650
<< psubdiffcont >>
rect 70 650 130 750
<< locali >>
rect 70 750 130 766
rect 70 634 130 650
<< viali >>
rect 80 660 120 740
<< metal1 >>
rect -200 1070 150 1110
rect -300 720 -240 1040
rect -200 910 -40 980
rect 200 910 260 1140
rect -200 850 260 910
rect -200 780 -40 850
rect 70 740 130 760
rect 70 690 80 740
rect -200 660 80 690
rect 120 690 130 740
rect 200 720 260 850
rect 480 780 620 1180
rect 120 660 650 690
rect -200 650 650 660
use sky130_fd_pr__nfet_01v8_9CME3F  XM1
timestamp 1665779562
transform 0 -1 -152 1 0 753
box -73 -148 73 148
use sky130_fd_pr__nfet_01v8_Z2KCLS  XM3
timestamp 1665882771
transform 0 -1 439 1 0 753
box -73 -239 73 239
use sky130_fd_pr__pfet_01v8_5AWN3K  sky130_fd_pr__pfet_01v8_5AWN3K_0
timestamp 1665779562
transform 0 -1 -71 1 0 1009
box -109 -263 109 229
use sky130_fd_pr__pfet_01v8_S6MTYS  sky130_fd_pr__pfet_01v8_S6MTYS_0
timestamp 1665882771
transform 0 -1 465 1 0 1061
box -161 -265 161 265
<< labels >>
rlabel metal1 -300 720 -240 1040 1 Vin
port 2 n
rlabel metal1 -200 650 650 690 1 VSS
port 4 n
<< end >>
