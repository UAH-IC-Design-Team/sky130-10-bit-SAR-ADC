magic
tech sky130A
magscale 1 2
timestamp 1666290788
<< metal3 >>
rect -1398 792 -626 820
rect -1398 368 -710 792
rect -646 368 -626 792
rect -1398 340 -626 368
rect -386 792 386 820
rect -386 368 302 792
rect 366 368 386 792
rect -386 340 386 368
rect 626 792 1398 820
rect 626 368 1314 792
rect 1378 368 1398 792
rect 626 340 1398 368
rect -1398 212 -626 240
rect -1398 -212 -710 212
rect -646 -212 -626 212
rect -1398 -240 -626 -212
rect -386 212 386 240
rect -386 -212 302 212
rect 366 -212 386 212
rect -386 -240 386 -212
rect 626 212 1398 240
rect 626 -212 1314 212
rect 1378 -212 1398 212
rect 626 -240 1398 -212
rect -1398 -368 -626 -340
rect -1398 -792 -710 -368
rect -646 -792 -626 -368
rect -1398 -820 -626 -792
rect -386 -368 386 -340
rect -386 -792 302 -368
rect 366 -792 386 -368
rect -386 -820 386 -792
rect 626 -368 1398 -340
rect 626 -792 1314 -368
rect 1378 -792 1398 -368
rect 626 -820 1398 -792
<< via3 >>
rect -710 368 -646 792
rect 302 368 366 792
rect 1314 368 1378 792
rect -710 -212 -646 212
rect 302 -212 366 212
rect 1314 -212 1378 212
rect -710 -792 -646 -368
rect 302 -792 366 -368
rect 1314 -792 1378 -368
<< mimcap >>
rect -1358 740 -958 780
rect -1358 420 -1318 740
rect -998 420 -958 740
rect -1358 380 -958 420
rect -346 740 54 780
rect -346 420 -306 740
rect 14 420 54 740
rect -346 380 54 420
rect 666 740 1066 780
rect 666 420 706 740
rect 1026 420 1066 740
rect 666 380 1066 420
rect -1358 160 -958 200
rect -1358 -160 -1318 160
rect -998 -160 -958 160
rect -1358 -200 -958 -160
rect -346 160 54 200
rect -346 -160 -306 160
rect 14 -160 54 160
rect -346 -200 54 -160
rect 666 160 1066 200
rect 666 -160 706 160
rect 1026 -160 1066 160
rect 666 -200 1066 -160
rect -1358 -420 -958 -380
rect -1358 -740 -1318 -420
rect -998 -740 -958 -420
rect -1358 -780 -958 -740
rect -346 -420 54 -380
rect -346 -740 -306 -420
rect 14 -740 54 -420
rect -346 -780 54 -740
rect 666 -420 1066 -380
rect 666 -740 706 -420
rect 1026 -740 1066 -420
rect 666 -780 1066 -740
<< mimcapcontact >>
rect -1318 420 -998 740
rect -306 420 14 740
rect 706 420 1026 740
rect -1318 -160 -998 160
rect -306 -160 14 160
rect 706 -160 1026 160
rect -1318 -740 -998 -420
rect -306 -740 14 -420
rect 706 -740 1026 -420
<< metal4 >>
rect -1210 741 -1106 870
rect -730 792 -626 870
rect -1319 740 -997 741
rect -1319 420 -1318 740
rect -998 420 -997 740
rect -1319 419 -997 420
rect -1210 161 -1106 419
rect -730 368 -710 792
rect -646 368 -626 792
rect -198 741 -94 870
rect 282 792 386 870
rect -307 740 15 741
rect -307 420 -306 740
rect 14 420 15 740
rect -307 419 15 420
rect -730 212 -626 368
rect -1319 160 -997 161
rect -1319 -160 -1318 160
rect -998 -160 -997 160
rect -1319 -161 -997 -160
rect -1210 -419 -1106 -161
rect -730 -212 -710 212
rect -646 -212 -626 212
rect -198 161 -94 419
rect 282 368 302 792
rect 366 368 386 792
rect 814 741 918 870
rect 1294 792 1398 870
rect 705 740 1027 741
rect 705 420 706 740
rect 1026 420 1027 740
rect 705 419 1027 420
rect 282 212 386 368
rect -307 160 15 161
rect -307 -160 -306 160
rect 14 -160 15 160
rect -307 -161 15 -160
rect -730 -368 -626 -212
rect -1319 -420 -997 -419
rect -1319 -740 -1318 -420
rect -998 -740 -997 -420
rect -1319 -741 -997 -740
rect -1210 -870 -1106 -741
rect -730 -792 -710 -368
rect -646 -792 -626 -368
rect -198 -419 -94 -161
rect 282 -212 302 212
rect 366 -212 386 212
rect 814 161 918 419
rect 1294 368 1314 792
rect 1378 368 1398 792
rect 1294 212 1398 368
rect 705 160 1027 161
rect 705 -160 706 160
rect 1026 -160 1027 160
rect 705 -161 1027 -160
rect 282 -368 386 -212
rect -307 -420 15 -419
rect -307 -740 -306 -420
rect 14 -740 15 -420
rect -307 -741 15 -740
rect -730 -870 -626 -792
rect -198 -870 -94 -741
rect 282 -792 302 -368
rect 366 -792 386 -368
rect 814 -419 918 -161
rect 1294 -212 1314 212
rect 1378 -212 1398 212
rect 1294 -368 1398 -212
rect 705 -420 1027 -419
rect 705 -740 706 -420
rect 1026 -740 1027 -420
rect 705 -741 1027 -740
rect 282 -870 386 -792
rect 814 -870 918 -741
rect 1294 -792 1314 -368
rect 1378 -792 1398 -368
rect 1294 -870 1398 -792
<< properties >>
string FIXED_BBOX 626 340 1106 820
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
