** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/controller/controller.sch
.subckt controller clk sw_n_sp9 sw_n_sp8 sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2
+ sw_n_sp1 VSS VDD reset sw_n8 sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6
+ sw_p_sp5 sw_p_sp4 sw_p_sp3 sw_p_sp2 sw_p_sp1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 bit10 bit9 bit8
+ bit7 bit6 bit5 bit4 bit3 bit2 bit1 done sw_sample comparator_clk comp_out_p comp_out_n
*.PININFO clk:I sw_n_sp[9..1]:O VSS:B VDD:B reset:I sw_n[8..1]:O sw_p_sp[9..1]:O sw_p[8..1]:O
*+ bit[10..1]:O done:O sw_sample:O comparator_clk:O comp_out_p:I comp_out_n:I
x3 VDD raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7 raw_bit6 raw_bit5 raw_bit4
+ raw_bit3 raw_bit2 raw_bit1 VSS reset bit10 bit9 bit8 bit7 bit6 bit5 bit4 bit3 bit2 bit1 done cycle13 dec
x4 raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7 raw_bit6 raw_bit5 raw_bit4
+ raw_bit3 raw_bit2 raw_bit1 cycle12 cycle11 cycle10 cycle9 cycle8 cycle7 cycle6 cycle5 cycle4 cycle3 cycle2
+ cycle1 cycle0 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 Vcmp_buff raw_bit_calc_reset VDD VSS
+ sw_n_sp9 sw_n_sp8 sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2 sw_n_sp1 sw_n8 sw_n7 sw_n6 sw_n5
+ sw_n4 sw_n3 sw_n2 sw_n1 sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6 sw_p_sp5 sw_p_sp4 sw_p_sp3 sw_p_sp2 sw_p_sp1
+ raw_bit_calculator
x1 VDD controller_clk sw_sample VSS reset cycle15 cycle14 cycle13 cycle12 cycle11 cycle10 cycle9
+ cycle8 cycle7 cycle6 cycle5 cycle4 cycle3 cycle2 cycle1 cycle0 shifted_clock_generator
x2 net1 reset VSS VSS VDD VDD net6 sky130_fd_sc_hd__and2_1
x6 cycle14 cycle15 VSS VSS VDD VDD net1 sky130_fd_sc_hd__xnor2_1
x25 net3 VSS VSS VDD VDD Vcmp_buff sky130_fd_sc_hd__buf_16
x26 comp_out_p VSS VSS VDD VDD net2 sky130_fd_sc_hd__buf_4
x27 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__buf_8
x28 net4 VSS VSS VDD VDD raw_bit_calc_reset sky130_fd_sc_hd__buf_16
x29 net6 VSS VSS VDD VDD net5 sky130_fd_sc_hd__buf_4
x30 net5 VSS VSS VDD VDD net4 sky130_fd_sc_hd__buf_8
x5 VDD clk reset VSS sw_sample comparator_clk sample_clock
x7 VSS comp_out_p VDD comp_out_n controller_clk xor_clock_gen
.ends

* expanding   symbol:  src/dec/dec.sym # of pins=7
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/dec/dec.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/dec/dec.sch
.subckt dec VDD raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7 raw_bit6 raw_bit5
+ raw_bit4 raw_bit3 raw_bit2 raw_bit1 VSS reset_b bit10 bit9 bit8 bit7 bit6 bit5 bit4 bit3 bit2 bit1 done
+ dump_bus
*.PININFO VDD:B bit[10..1]:O VSS:B reset_b:I dump_bus:I done:O raw_bit[13..1]:I
x62 raw_bit2 raw_bit1 net1 VSS VSS VDD VDD net16 net2 sky130_fd_sc_hd__fa_1
x64 raw_bit3 raw_bit1 net4 VSS VSS VDD VDD net1 net3 sky130_fd_sc_hd__fa_1
x67 dump_bus net2 reset_b VSS VSS VDD VDD bit2 sky130_fd_sc_hd__dfrtp_1
x68 dump_bus net3 reset_b VSS VSS VDD VDD bit3 sky130_fd_sc_hd__dfrtp_1
x65 raw_bit5 raw_bit4 net5 VSS VSS VDD VDD net4 net6 sky130_fd_sc_hd__fa_1
x69 raw_bit6 raw_bit4 net8 VSS VSS VDD VDD net5 net7 sky130_fd_sc_hd__fa_1
x70 dump_bus net6 reset_b VSS VSS VDD VDD bit4 sky130_fd_sc_hd__dfrtp_1
x71 dump_bus net7 reset_b VSS VSS VDD VDD bit5 sky130_fd_sc_hd__dfrtp_1
x72 raw_bit7 raw_bit4 net9 VSS VSS VDD VDD net8 net10 sky130_fd_sc_hd__fa_1
x73 raw_bit9 raw_bit8 net12 VSS VSS VDD VDD net9 net11 sky130_fd_sc_hd__fa_1
x74 dump_bus net10 reset_b VSS VSS VDD VDD bit6 sky130_fd_sc_hd__dfrtp_1
x75 dump_bus net11 reset_b VSS VSS VDD VDD bit7 sky130_fd_sc_hd__dfrtp_1
x76 raw_bit10 raw_bit8 net13 VSS VSS VDD VDD net12 net14 sky130_fd_sc_hd__fa_1
x77 raw_bit11 raw_bit8 raw_bit12 VSS VSS VDD VDD net13 net15 sky130_fd_sc_hd__fa_1
x78 dump_bus net14 reset_b VSS VSS VDD VDD bit8 sky130_fd_sc_hd__dfrtp_1
x79 dump_bus net15 reset_b VSS VSS VDD VDD bit9 sky130_fd_sc_hd__dfrtp_1
x80 dump_bus net16 reset_b VSS VSS VDD VDD bit1 sky130_fd_sc_hd__dfrtp_1
x81 dump_bus raw_bit13 reset_b VSS VSS VDD VDD bit10 sky130_fd_sc_hd__dfrtp_1
x82 dump_bus VSS VSS VDD VDD done sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  src/raw_bit_calculator/raw_bit_calculator.sym # of pins=10
** sym_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/raw_bit_calculator/raw_bit_calculator.sym
** sch_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/raw_bit_calculator/raw_bit_calculator.sch
.subckt raw_bit_calculator raw_bit13 raw_bit12 raw_bit11 raw_bit10 raw_bit9 raw_bit8 raw_bit7
+ raw_bit6 raw_bit5 raw_bit4 raw_bit3 raw_bit2 raw_bit1 cycle13 cycle12 cycle11 cycle10 cycle9 cycle8 cycle7
+ cycle6 cycle5 cycle4 cycle3 cycle2 cycle1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 Vcmp RESET VDD
+ VSS sw_n_sp9 sw_n_sp8 sw_n_sp7 sw_n_sp6 sw_n_sp5 sw_n_sp4 sw_n_sp3 sw_n_sp2 sw_n_sp1 sw_n8 sw_n7 sw_n6
+ sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 sw_p_sp9 sw_p_sp8 sw_p_sp7 sw_p_sp6 sw_p_sp5 sw_p_sp4 sw_p_sp3 sw_p_sp2
+ sw_p_sp1
*.PININFO cycle[13..1]:I sw_n_sp[9..1]:O VSS:B VDD:B sw_n[8..1]:O sw_p_sp[9..1]:O sw_p[8..1]:O
*+ Vcmp:I RESET:I raw_bit[13..1]:O
x29 raw_bit1 Vcmp VSS VSS VDD VDD net58 sky130_fd_sc_hd__xor2_1
x31 raw_bit1 Vcmp VSS VSS VDD VDD net62 sky130_fd_sc_hd__xor2_1
x37 raw_bit4 Vcmp VSS VSS VDD VDD net52 sky130_fd_sc_hd__xor2_1
x40 raw_bit4 Vcmp VSS VSS VDD VDD net53 sky130_fd_sc_hd__xor2_1
x45 raw_bit4 Vcmp VSS VSS VDD VDD net54 sky130_fd_sc_hd__xor2_1
x100 cycle1 net11 net23 VSS VSS VDD VDD sw_p_sp1 sky130_fd_sc_hd__dfrtp_1
x99 Vcmp VSS VSS VDD VDD net11 sky130_fd_sc_hd__inv_1
x102 cycle1 Vcmp net23 VSS VSS VDD VDD sw_n_sp1 sky130_fd_sc_hd__dfrtp_1
x25 cycle1 Vcmp net25 VSS VSS VDD VDD sw_n_sp2 sky130_fd_sc_hd__dfrtp_1
x103 Vcmp VSS VSS VDD VDD net12 sky130_fd_sc_hd__inv_1
x104 cycle1 net12 net25 VSS VSS VDD VDD sw_p_sp2 sky130_fd_sc_hd__dfrtp_1
x21 net1 Vcmp RESET VSS VSS VDD VDD sw_n1 sky130_fd_sc_hd__dfstp_1
x22 net1 net13 RESET VSS VSS VDD VDD sw_p1 sky130_fd_sc_hd__dfstp_1
x105 Vcmp VSS VSS VDD VDD net13 sky130_fd_sc_hd__inv_1
x28 net4 Vcmp RESET VSS VSS VDD VDD sw_n2 sky130_fd_sc_hd__dfstp_1
x106 net4 net14 RESET VSS VSS VDD VDD sw_p2 sky130_fd_sc_hd__dfstp_1
x107 Vcmp VSS VSS VDD VDD net14 sky130_fd_sc_hd__inv_1
x109 Vcmp VSS VSS VDD VDD net15 sky130_fd_sc_hd__inv_1
x111 Vcmp VSS VSS VDD VDD net16 sky130_fd_sc_hd__inv_1
x27 cycle4 Vcmp net27 VSS VSS VDD VDD sw_n_sp3 sky130_fd_sc_hd__dfrtp_1
x35 cycle4 net15 net27 VSS VSS VDD VDD sw_p_sp3 sky130_fd_sc_hd__dfrtp_1
x41 cycle4 Vcmp net28 VSS VSS VDD VDD sw_n_sp4 sky130_fd_sc_hd__dfrtp_1
x108 cycle4 net16 net28 VSS VSS VDD VDD sw_p_sp4 sky130_fd_sc_hd__dfrtp_1
x110 cycle4 Vcmp net29 VSS VSS VDD VDD sw_n_sp5 sky130_fd_sc_hd__dfrtp_1
x112 cycle4 net17 net29 VSS VSS VDD VDD sw_p_sp5 sky130_fd_sc_hd__dfrtp_1
x113 Vcmp VSS VSS VDD VDD net17 sky130_fd_sc_hd__inv_1
x114 net6 net18 RESET VSS VSS VDD VDD sw_p3 sky130_fd_sc_hd__dfstp_1
x32 net6 Vcmp RESET VSS VSS VDD VDD sw_n3 sky130_fd_sc_hd__dfstp_1
x115 Vcmp VSS VSS VDD VDD net18 sky130_fd_sc_hd__inv_1
x38 net7 Vcmp RESET VSS VSS VDD VDD sw_n4 sky130_fd_sc_hd__dfstp_1
x116 net7 net19 RESET VSS VSS VDD VDD sw_p4 sky130_fd_sc_hd__dfstp_1
x117 Vcmp VSS VSS VDD VDD net19 sky130_fd_sc_hd__inv_1
x43 net8 Vcmp RESET VSS VSS VDD VDD sw_n5 sky130_fd_sc_hd__dfstp_1
x118 net8 net20 RESET VSS VSS VDD VDD sw_p5 sky130_fd_sc_hd__dfstp_1
x119 Vcmp VSS VSS VDD VDD net20 sky130_fd_sc_hd__inv_1
x132 cycle12 net21 RESET VSS VSS VDD VDD sw_p_sp9 sky130_fd_sc_hd__dfrtp_1
x133 Vcmp VSS VSS VDD VDD net21 sky130_fd_sc_hd__inv_1
x61 cycle12 Vcmp RESET VSS VSS VDD VDD sw_n_sp9 sky130_fd_sc_hd__dfrtp_1
x24 net51 VDD VSS net1 net3 net2 demux2
x30 net61 VDD VSS net4 net60 net5 demux2
x34 net65 VDD VSS net6 net64 net22 demux2
x39 net68 VDD VSS net7 net67 net9 demux2
x44 net71 VDD VSS net8 net70 net10 demux2
x1 net2 VSS VSS VDD VDD net24 sky130_fd_sc_hd__inv_1
x2 net5 VSS VSS VDD VDD net26 sky130_fd_sc_hd__inv_1
x3 cycle1 Vcmp RESET VSS VSS VDD VDD raw_bit1 sky130_fd_sc_hd__dfrtp_4
x4 cycle2 Vcmp RESET VSS VSS VDD VDD raw_bit2 sky130_fd_sc_hd__dfrtp_4
x5 cycle3 Vcmp RESET VSS VSS VDD VDD raw_bit3 sky130_fd_sc_hd__dfrtp_4
x6 cycle4 Vcmp RESET VSS VSS VDD VDD raw_bit4 sky130_fd_sc_hd__dfrtp_4
x7 cycle5 Vcmp RESET VSS VSS VDD VDD raw_bit5 sky130_fd_sc_hd__dfrtp_4
x8 cycle6 Vcmp RESET VSS VSS VDD VDD raw_bit6 sky130_fd_sc_hd__dfrtp_4
x9 cycle7 Vcmp RESET VSS VSS VDD VDD raw_bit7 sky130_fd_sc_hd__dfrtp_4
x10 cycle8 Vcmp RESET VSS VSS VDD VDD raw_bit8 sky130_fd_sc_hd__dfrtp_4
x11 cycle9 Vcmp RESET VSS VSS VDD VDD raw_bit9 sky130_fd_sc_hd__dfrtp_4
x12 cycle10 Vcmp RESET VSS VSS VDD VDD raw_bit10 sky130_fd_sc_hd__dfrtp_4
x13 cycle11 Vcmp RESET VSS VSS VDD VDD raw_bit11 sky130_fd_sc_hd__dfrtp_4
x14 cycle12 Vcmp RESET VSS VSS VDD VDD raw_bit12 sky130_fd_sc_hd__dfrtp_4
x15 cycle13 Vcmp RESET VSS VSS VDD VDD raw_bit13 sky130_fd_sc_hd__dfrtp_4
x18 net22 VSS VSS VDD VDD net30 sky130_fd_sc_hd__inv_1
x19 net9 VSS VSS VDD VDD net31 sky130_fd_sc_hd__inv_1
x20 net10 VSS VSS VDD VDD net32 sky130_fd_sc_hd__inv_1
x42 raw_bit8 Vcmp VSS VSS VDD VDD net55 sky130_fd_sc_hd__xor2_1
x62 raw_bit8 Vcmp VSS VSS VDD VDD net56 sky130_fd_sc_hd__xor2_1
x64 raw_bit8 Vcmp VSS VSS VDD VDD net57 sky130_fd_sc_hd__xor2_1
x65 Vcmp VSS VSS VDD VDD net38 sky130_fd_sc_hd__inv_1
x66 Vcmp VSS VSS VDD VDD net39 sky130_fd_sc_hd__inv_1
x67 cycle8 Vcmp net45 VSS VSS VDD VDD sw_n_sp6 sky130_fd_sc_hd__dfrtp_1
x68 cycle8 net38 net45 VSS VSS VDD VDD sw_p_sp6 sky130_fd_sc_hd__dfrtp_1
x69 cycle8 Vcmp net46 VSS VSS VDD VDD sw_n_sp7 sky130_fd_sc_hd__dfrtp_1
x70 cycle8 net39 net46 VSS VSS VDD VDD sw_p_sp7 sky130_fd_sc_hd__dfrtp_1
x71 cycle8 Vcmp net47 VSS VSS VDD VDD sw_n_sp8 sky130_fd_sc_hd__dfrtp_1
x72 cycle8 net40 net47 VSS VSS VDD VDD sw_p_sp8 sky130_fd_sc_hd__dfrtp_1
x73 Vcmp VSS VSS VDD VDD net40 sky130_fd_sc_hd__inv_1
x74 net33 net41 RESET VSS VSS VDD VDD sw_p6 sky130_fd_sc_hd__dfstp_1
x75 net33 Vcmp RESET VSS VSS VDD VDD sw_n6 sky130_fd_sc_hd__dfstp_1
x76 Vcmp VSS VSS VDD VDD net41 sky130_fd_sc_hd__inv_1
x77 net34 Vcmp RESET VSS VSS VDD VDD sw_n7 sky130_fd_sc_hd__dfstp_1
x78 net34 net42 RESET VSS VSS VDD VDD sw_p7 sky130_fd_sc_hd__dfstp_1
x79 Vcmp VSS VSS VDD VDD net42 sky130_fd_sc_hd__inv_1
x80 net35 Vcmp RESET VSS VSS VDD VDD sw_n8 sky130_fd_sc_hd__dfstp_1
x81 net35 net43 RESET VSS VSS VDD VDD sw_p8 sky130_fd_sc_hd__dfstp_1
x82 Vcmp VSS VSS VDD VDD net43 sky130_fd_sc_hd__inv_1
x83 net74 VDD VSS net33 net73 net44 demux2
x84 net77 VDD VSS net34 net76 net36 demux2
x85 net80 VDD VSS net35 net79 net37 demux2
x88 net44 VSS VSS VDD VDD net48 sky130_fd_sc_hd__inv_1
x89 net36 VSS VSS VDD VDD net49 sky130_fd_sc_hd__inv_1
x90 net37 VSS VSS VDD VDD net50 sky130_fd_sc_hd__inv_1
x46 net24 RESET VSS VSS VDD VDD net23 sky130_fd_sc_hd__and2_0
x23 net26 RESET VSS VSS VDD VDD net25 sky130_fd_sc_hd__and2_0
x26 net30 RESET VSS VSS VDD VDD net27 sky130_fd_sc_hd__and2_0
x16 net31 RESET VSS VSS VDD VDD net28 sky130_fd_sc_hd__and2_0
x17 net32 RESET VSS VSS VDD VDD net29 sky130_fd_sc_hd__and2_0
x33 net48 RESET VSS VSS VDD VDD net45 sky130_fd_sc_hd__and2_0
x36 net49 RESET VSS VSS VDD VDD net46 sky130_fd_sc_hd__and2_0
x47 net50 RESET VSS VSS VDD VDD net47 sky130_fd_sc_hd__and2_0
x48 cycle2 net58 RESET VSS VSS VDD VDD net51 sky130_fd_sc_hd__dfrtp_1
x49 net59 VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkdlybuf4s50_1
x50 cycle2 VSS VSS VDD VDD net59 sky130_fd_sc_hd__clkdlybuf4s50_1
x51 cycle3 net62 RESET VSS VSS VDD VDD net61 sky130_fd_sc_hd__dfrtp_1
x52 net63 VSS VSS VDD VDD net60 sky130_fd_sc_hd__clkdlybuf4s50_1
x53 cycle3 VSS VSS VDD VDD net63 sky130_fd_sc_hd__clkdlybuf4s50_1
x54 cycle5 net52 RESET VSS VSS VDD VDD net65 sky130_fd_sc_hd__dfrtp_1
x55 net66 VSS VSS VDD VDD net64 sky130_fd_sc_hd__clkdlybuf4s50_1
x56 cycle5 VSS VSS VDD VDD net66 sky130_fd_sc_hd__clkdlybuf4s50_1
x57 cycle6 net53 RESET VSS VSS VDD VDD net68 sky130_fd_sc_hd__dfrtp_1
x58 net69 VSS VSS VDD VDD net67 sky130_fd_sc_hd__clkdlybuf4s50_1
x59 cycle6 VSS VSS VDD VDD net69 sky130_fd_sc_hd__clkdlybuf4s50_1
x60 cycle7 net54 RESET VSS VSS VDD VDD net71 sky130_fd_sc_hd__dfrtp_1
x63 net72 VSS VSS VDD VDD net70 sky130_fd_sc_hd__clkdlybuf4s50_1
x86 cycle7 VSS VSS VDD VDD net72 sky130_fd_sc_hd__clkdlybuf4s50_1
x87 cycle9 net55 RESET VSS VSS VDD VDD net74 sky130_fd_sc_hd__dfrtp_1
x91 net75 VSS VSS VDD VDD net73 sky130_fd_sc_hd__clkdlybuf4s50_1
x92 cycle9 VSS VSS VDD VDD net75 sky130_fd_sc_hd__clkdlybuf4s50_1
x93 cycle10 net56 RESET VSS VSS VDD VDD net77 sky130_fd_sc_hd__dfrtp_1
x94 net78 VSS VSS VDD VDD net76 sky130_fd_sc_hd__clkdlybuf4s50_1
x95 cycle10 VSS VSS VDD VDD net78 sky130_fd_sc_hd__clkdlybuf4s50_1
x96 cycle11 net57 RESET VSS VSS VDD VDD net80 sky130_fd_sc_hd__dfrtp_1
x97 net81 VSS VSS VDD VDD net79 sky130_fd_sc_hd__clkdlybuf4s50_1
x98 cycle11 VSS VSS VDD VDD net81 sky130_fd_sc_hd__clkdlybuf4s50_1
.ends


* expanding   symbol:  src/shifted_clock_generator/shifted_clock_generator.sym # of pins=6
** sym_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/shifted_clock_generator/shifted_clock_generator.sym
** sch_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/shifted_clock_generator/shifted_clock_generator.sch
.subckt shifted_clock_generator VDD clk sw_sample VSS reset cycle15 cycle14 cycle13 cycle12 cycle11
+ cycle10 cycle9 cycle8 cycle7 cycle6 cycle5 cycle4 cycle3 cycle2 cycle1 cycle0
*.PININFO cycle[15..0]:O VSS:B VDD:B clk:I reset:I sw_sample:I
x32 net16 net17 reset_b VSS VSS VDD VDD net4 sky130_fd_sc_hd__dfrtp_1
x1 net5 net4 reset_b VSS VSS VDD VDD net18 sky130_fd_sc_hd__dfrtp_1
x2 net6 net18 reset_b VSS VSS VDD VDD net19 sky130_fd_sc_hd__dfrtp_1
x3 net7 net19 reset_b VSS VSS VDD VDD net20 sky130_fd_sc_hd__dfrtp_1
x4 net8 net20 reset_b VSS VSS VDD VDD net21 sky130_fd_sc_hd__dfrtp_1
x5 net9 net21 reset_b VSS VSS VDD VDD net22 sky130_fd_sc_hd__dfrtp_1
x6 net10 net22 reset_b VSS VSS VDD VDD net23 sky130_fd_sc_hd__dfrtp_1
x7 net11 net23 reset_b VSS VSS VDD VDD net24 sky130_fd_sc_hd__dfrtp_1
x8 net12 net24 reset_b VSS VSS VDD VDD net25 sky130_fd_sc_hd__dfrtp_1
x9 net13 net25 reset_b VSS VSS VDD VDD net26 sky130_fd_sc_hd__dfrtp_1
x10 net14 net26 reset_b VSS VSS VDD VDD net27 sky130_fd_sc_hd__dfrtp_1
x11 net15 net27 reset_b VSS VSS VDD VDD net28 sky130_fd_sc_hd__dfrtp_1
x12 net3 net28 reset_b VSS VSS VDD VDD net29 sky130_fd_sc_hd__dfrtp_1
x13 net1 net29 reset_b VSS VSS VDD VDD net30 sky130_fd_sc_hd__dfrtp_1
x14 net2 net30 reset_b VSS VSS VDD VDD net31 sky130_fd_sc_hd__dfrtp_1
x31 net32 net33 reset_b VSS VSS VDD VDD net17 sky130_fd_sc_hd__dfrtp_1
x37 net35 VSS VSS VDD VDD reset_b sky130_fd_sc_hd__buf_16
x35 net34 reset VSS VSS VDD VDD net35 sky130_fd_sc_hd__and2_4
x15 net17 VSS VSS VDD VDD net46 sky130_fd_sc_hd__buf_1
x16 net44 VSS VSS VDD VDD net36 sky130_fd_sc_hd__buf_2
x20 net44 VSS VSS VDD VDD net37 sky130_fd_sc_hd__buf_2
x21 net44 VSS VSS VDD VDD net38 sky130_fd_sc_hd__buf_2
x22 net44 VSS VSS VDD VDD net39 sky130_fd_sc_hd__buf_2
x23 net45 VSS VSS VDD VDD net40 sky130_fd_sc_hd__buf_2
x24 net45 VSS VSS VDD VDD net41 sky130_fd_sc_hd__buf_2
x25 net45 VSS VSS VDD VDD net42 sky130_fd_sc_hd__buf_2
x26 net45 VSS VSS VDD VDD net43 sky130_fd_sc_hd__buf_2
x27 clk VSS VSS VDD VDD net44 sky130_fd_sc_hd__buf_4
x28 clk VSS VSS VDD VDD net45 sky130_fd_sc_hd__buf_4
x17 net36 VSS VSS VDD VDD net32 sky130_fd_sc_hd__buf_1
x18 net36 VSS VSS VDD VDD net16 sky130_fd_sc_hd__buf_1
x19 net37 VSS VSS VDD VDD net5 sky130_fd_sc_hd__buf_1
x29 net37 VSS VSS VDD VDD net6 sky130_fd_sc_hd__buf_1
x30 net38 VSS VSS VDD VDD net7 sky130_fd_sc_hd__buf_1
x33 net38 VSS VSS VDD VDD net8 sky130_fd_sc_hd__buf_1
x47 net39 VSS VSS VDD VDD net9 sky130_fd_sc_hd__buf_1
x48 net39 VSS VSS VDD VDD net10 sky130_fd_sc_hd__buf_1
x51 net40 VSS VSS VDD VDD net11 sky130_fd_sc_hd__buf_1
x52 net40 VSS VSS VDD VDD net12 sky130_fd_sc_hd__buf_1
x53 net41 VSS VSS VDD VDD net13 sky130_fd_sc_hd__buf_1
x54 net41 VSS VSS VDD VDD net14 sky130_fd_sc_hd__buf_1
x55 net42 VSS VSS VDD VDD net15 sky130_fd_sc_hd__buf_1
x56 net42 VSS VSS VDD VDD net3 sky130_fd_sc_hd__buf_1
x57 net43 VSS VSS VDD VDD net1 sky130_fd_sc_hd__buf_1
x58 net43 VSS VSS VDD VDD net2 sky130_fd_sc_hd__buf_1
x62 net4 VSS VSS VDD VDD net47 sky130_fd_sc_hd__buf_1
x66 net18 VSS VSS VDD VDD net48 sky130_fd_sc_hd__buf_1
x70 net19 VSS VSS VDD VDD net49 sky130_fd_sc_hd__buf_1
x34 sw_sample VSS VSS VDD VDD net34 sky130_fd_sc_hd__inv_1
x36 VDD VSS VSS VDD VDD net33 sky130_fd_sc_hd__buf_1
x38 net46 VSS VSS VDD VDD cycle0 sky130_fd_sc_hd__buf_4
x39 net47 VSS VSS VDD VDD cycle1 sky130_fd_sc_hd__buf_4
x40 net48 VSS VSS VDD VDD cycle2 sky130_fd_sc_hd__buf_4
x41 net49 VSS VSS VDD VDD cycle3 sky130_fd_sc_hd__buf_4
x42 net20 VSS VSS VDD VDD net50 sky130_fd_sc_hd__buf_1
x43 net21 VSS VSS VDD VDD net51 sky130_fd_sc_hd__buf_1
x44 net22 VSS VSS VDD VDD net52 sky130_fd_sc_hd__buf_1
x45 net23 VSS VSS VDD VDD net53 sky130_fd_sc_hd__buf_1
x46 net50 VSS VSS VDD VDD cycle4 sky130_fd_sc_hd__buf_4
x49 net51 VSS VSS VDD VDD cycle5 sky130_fd_sc_hd__buf_4
x50 net52 VSS VSS VDD VDD cycle6 sky130_fd_sc_hd__buf_4
x59 net53 VSS VSS VDD VDD cycle7 sky130_fd_sc_hd__buf_4
x60 net24 VSS VSS VDD VDD net54 sky130_fd_sc_hd__buf_1
x61 net25 VSS VSS VDD VDD net55 sky130_fd_sc_hd__buf_1
x63 net26 VSS VSS VDD VDD net56 sky130_fd_sc_hd__buf_1
x64 net27 VSS VSS VDD VDD net57 sky130_fd_sc_hd__buf_1
x65 net54 VSS VSS VDD VDD cycle8 sky130_fd_sc_hd__buf_4
x67 net55 VSS VSS VDD VDD cycle9 sky130_fd_sc_hd__buf_4
x68 net56 VSS VSS VDD VDD cycle10 sky130_fd_sc_hd__buf_4
x69 net57 VSS VSS VDD VDD cycle11 sky130_fd_sc_hd__buf_4
x71 net28 VSS VSS VDD VDD net58 sky130_fd_sc_hd__buf_1
x72 net29 VSS VSS VDD VDD net59 sky130_fd_sc_hd__buf_1
x73 net30 VSS VSS VDD VDD net60 sky130_fd_sc_hd__buf_1
x74 net31 VSS VSS VDD VDD net61 sky130_fd_sc_hd__buf_1
x75 net58 VSS VSS VDD VDD cycle12 sky130_fd_sc_hd__buf_4
x76 net59 VSS VSS VDD VDD cycle13 sky130_fd_sc_hd__buf_4
x77 net60 VSS VSS VDD VDD cycle14 sky130_fd_sc_hd__buf_4
x78 net61 VSS VSS VDD VDD cycle15 sky130_fd_sc_hd__buf_4
.ends


* expanding   symbol:  src/sample_clock/sample_clock.sym # of pins=6
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/sample_clock/sample_clock.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/sample_clock/sample_clock.sch
.subckt sample_clock VDD clk reset VSS sw_sample comparator_clk
*.PININFO VDD:B clk:I sw_sample:O VSS:B comparator_clk:O reset:I
x5 clk johnson_counter_loop reset VSS VSS VDD VDD net1 sky130_fd_sc_hd__dfrtp_1
x7 clk net1 reset VSS VSS VDD VDD net2 sky130_fd_sc_hd__dfrtp_1
x8 clk net2 reset VSS VSS VDD VDD net3 sky130_fd_sc_hd__dfrtp_1
x9 clk net3 reset VSS VSS VDD VDD net4 sky130_fd_sc_hd__dfrtp_1
x10 clk net4 reset VSS VSS VDD VDD net5 sky130_fd_sc_hd__dfrtp_1
x11 clk net5 reset VSS VSS VDD VDD net6 sky130_fd_sc_hd__dfrtp_1
x12 clk net6 reset VSS VSS VDD VDD net7 sky130_fd_sc_hd__dfrtp_1
x13 clk net7 reset VSS VSS VDD VDD some_net sky130_fd_sc_hd__dfrtp_1
x14 clk some_net reset VSS VSS VDD VDD net8 sky130_fd_sc_hd__dfrtp_1
x15 clk net8 reset VSS VSS VDD VDD net9 sky130_fd_sc_hd__dfrtp_1
x16 clk net9 reset VSS VSS VDD VDD net10 sky130_fd_sc_hd__dfrtp_1
x17 clk net10 reset VSS VSS VDD VDD net11 sky130_fd_sc_hd__dfrtp_1
x18 clk net11 reset VSS VSS VDD VDD net12 sky130_fd_sc_hd__dfrtp_1
x19 clk net12 reset VSS VSS VDD VDD net13 sky130_fd_sc_hd__dfrtp_1
x20 clk net13 reset VSS VSS VDD VDD net14 sky130_fd_sc_hd__dfrtp_1
x21 clk net14 reset VSS VSS VDD VDD net15 sky130_fd_sc_hd__dfrtp_1
x22 net15 VSS VSS VDD VDD johnson_counter_loop sky130_fd_sc_hd__inv_1
x23 net17 net16 VSS VSS VDD VDD net20 sky130_fd_sc_hd__and2_1
x24 sw_sample VSS VSS VDD VDD net16 sky130_fd_sc_hd__inv_1
x25 net19 VSS VSS VDD VDD comparator_clk sky130_fd_sc_hd__buf_16
x26 net21 VSS VSS VDD VDD net18 sky130_fd_sc_hd__buf_4
x27 net18 VSS VSS VDD VDD net19 sky130_fd_sc_hd__buf_8
x1 net20 VSS VSS VDD VDD net21 sky130_fd_sc_hd__buf_2
x2 net23 VSS VSS VDD VDD net22 sky130_fd_sc_hd__buf_4
x3 net22 VSS VSS VDD VDD sw_sample sky130_fd_sc_hd__buf_8
x4 net1 VSS VSS VDD VDD net23 sky130_fd_sc_hd__buf_2
x6 net24 VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkdlybuf4s50_1
x28 clk VSS VSS VDD VDD net24 sky130_fd_sc_hd__clkdlybuf4s50_1
.ends


* expanding   symbol:  src/xor_clock_gen/xor_clock_gen.sym # of pins=5
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/xor_clock_gen/xor_clock_gen.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/xor_clock_gen/xor_clock_gen.sch
.subckt xor_clock_gen VSS Vin_p VDD Vin_n Gen_clk
*.PININFO Vin_p:I VSS:B Gen_clk:O VDD:B Vin_n:I
x2 Vin_p Vin_n VSS VSS VDD VDD net1 sky130_fd_sc_hd__xor2_1
x3 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__clkdlybuf4s50_1
x17 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkdlybuf4s50_1
x9 net11 VSS VSS VDD VDD net4 sky130_fd_sc_hd__clkbuf_1
x14 net4 VSS VSS VDD VDD net5 sky130_fd_sc_hd__clkbuf_2
x19 net5 VSS VSS VDD VDD net6 sky130_fd_sc_hd__clkbuf_4
x26 net6 VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkbuf_8
x27 net7 VSS VSS VDD VDD Gen_clk sky130_fd_sc_hd__clkbuf_16
XC1 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=3 m=3
x1 net3 VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkdlybuf4s50_1
x4 net9 VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkdlybuf4s50_1
x5 net8 VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkdlybuf4s50_1
x6 net10 VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkdlybuf4s50_1
.ends


* expanding   symbol:  src/demux2/demux2.sym # of pins=6
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sch
.subckt demux2 S VDD VSS OUT_0 IN OUT_1
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
x1 net1 IN VSS VSS VDD VDD OUT_0 sky130_fd_sc_hd__and2_0
x2 S IN VSS VSS VDD VDD OUT_1 sky130_fd_sc_hd__and2_0
x3 S VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_1
.ends

.end
