** sch_path:
*+ /foss/designs/sky130-10-bit-SAR-ADC/xschem/tests/pulse_generator/pulse_generator_test.sch
**.subckt pulse_generator_test
V1 clk GND PULSE 0 1.8 20us 1ns 1ns 5us 10us
V2 RST_PLS GND PULSE 1.8V 0 0 1ns 1ns 5us 1s
x2 clk Pulse VDD VSS RST_PLS pulse_generator
V3 VDD GND 1.8V
V4 VSS GND 0
**** begin user architecture code
 .lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice



.options acct list
.temp 25
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
.control
tran 0.1u 400u
plot RST_PLS clk+2 Pulse+4
write pulse_generator_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  src/pulse_generator/pulse_generator.sym # of pins=5
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/pulse_generator/pulse_generator.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/pulse_generator/pulse_generator.sch
.subckt pulse_generator  clk pulse VDD VSS RST_PLS
*.ipin clk
*.ipin RST_PLS
*.opin pulse
*.iopin VDD
*.iopin VSS
x1 clk net1 RST_PLS VSS VSS VDD VDD clk2 net1 sky130_fd_sc_hd__dfrbp_1
x2 clk2 net2 RST_PLS VSS VSS VDD VDD clk4 net2 sky130_fd_sc_hd__dfrbp_1
x3 clk4 net3 RST_PLS VSS VSS VDD VDD clk8 net3 sky130_fd_sc_hd__dfrbp_1
x4 clk8 net4 RST_PLS VSS VSS VDD VDD clk16 net4 sky130_fd_sc_hd__dfrbp_1
x5 delayed clk64 VSS VSS VDD VDD net7 sky130_fd_sc_hd__xor2_1
x9 clk16 net5 RST_PLS VSS VSS VDD VDD clk32 net5 sky130_fd_sc_hd__dfrbp_1
x10 clk32 net6 RST_PLS VSS VSS VDD VDD clk64 net6 sky130_fd_sc_hd__dfrbp_1
x6 clk clk64 RST_PLS VSS VSS VDD VDD delayed sky130_fd_sc_hd__dfrtp_1
x7 clk net7 RST_PLS VSS VSS VDD VDD pulse sky130_fd_sc_hd__dfrtn_1
.ends

.GLOBAL GND
.end
