magic
tech sky130A
timestamp 1667663783
<< metal4 >>
rect 250 5200 310 5800
rect 590 5200 650 5800
rect 1050 5200 1110 5800
rect 1390 5200 1450 5800
rect 1850 5200 1910 5800
rect 2190 5200 2250 5800
rect 2650 5200 2710 5800
rect 2990 5200 3050 5800
rect 3450 5200 3510 5800
rect 3790 5200 3850 5800
rect 4250 5200 4310 5800
rect 4590 5200 4650 5800
rect 5050 5200 5110 5800
rect 5390 5200 5450 5800
rect 5850 5200 5910 5800
rect 6190 5200 6250 5800
rect 6650 5200 6710 5800
rect 6990 5200 7050 5800
rect 7450 5200 7510 5800
rect 7790 5200 7850 5800
rect 8250 5200 8310 5800
rect 8590 5200 8650 5800
rect 9050 5200 9110 5800
rect 9390 5200 9450 5800
rect 9850 5200 9910 5800
rect 10190 5200 10250 5800
rect 10650 5200 10710 5800
rect 10990 5200 11050 5800
rect 11450 5200 11510 5800
rect 11790 5200 11850 5800
rect 12250 5200 12310 5800
rect 12590 5200 12650 5800
rect 250 4400 310 5000
rect 590 4400 650 5000
rect 1050 4400 1110 5000
rect 1390 4400 1450 5000
rect 1850 4400 1910 5000
rect 2190 4400 2250 5000
rect 2650 4400 2710 5000
rect 2990 4400 3050 5000
rect 3450 4400 3510 5000
rect 3790 4400 3850 5000
rect 4250 4400 4310 5000
rect 4590 4400 4650 5000
rect 5050 4400 5110 5000
rect 5390 4400 5450 5000
rect 5850 4400 5910 5000
rect 6190 4400 6250 5000
rect 6650 4400 6710 5000
rect 6990 4400 7050 5000
rect 7450 4400 7510 5000
rect 7790 4400 7850 5000
rect 8250 4400 8310 5000
rect 8590 4400 8650 5000
rect 9050 4400 9110 5000
rect 9390 4400 9450 5000
rect 9850 4400 9910 5000
rect 10190 4400 10250 5000
rect 10650 4400 10710 5000
rect 10990 4400 11050 5000
rect 11450 4400 11510 5000
rect 11790 4400 11850 5000
rect 12250 4400 12310 5000
rect 12590 4400 12650 5000
rect 250 3600 310 4200
rect 590 3600 650 4200
rect 1050 3600 1110 4200
rect 1390 3600 1450 4200
rect 1850 3600 1910 4200
rect 2190 3600 2250 4200
rect 2650 3600 2710 4200
rect 2990 3600 3050 4200
rect 3450 3600 3510 4200
rect 3790 3600 3850 4200
rect 4250 3600 4310 4200
rect 4590 3600 4650 4200
rect 5050 3600 5110 4200
rect 5390 3600 5450 4200
rect 5850 3600 5910 4200
rect 6190 3600 6250 4200
rect 6650 3600 6710 4200
rect 6990 3600 7050 4200
rect 7450 3600 7510 4200
rect 7790 3600 7850 4200
rect 8250 3600 8310 4200
rect 8590 3600 8650 4200
rect 9050 3600 9110 4200
rect 9390 3600 9450 4200
rect 9850 3600 9910 4200
rect 10190 3600 10250 4200
rect 10650 3600 10710 4200
rect 10990 3600 11050 4200
rect 11450 3600 11510 4200
rect 11790 3600 11850 4200
rect 12250 3600 12310 4200
rect 12590 3600 12650 4200
rect 250 2800 310 3400
rect 590 2800 650 3400
rect 1050 2800 1110 3400
rect 1390 2800 1450 3400
rect 1850 2800 1910 3400
rect 2190 2800 2250 3400
rect 2650 2800 2710 3400
rect 2990 2800 3050 3400
rect 3450 2800 3510 3400
rect 3790 2800 3850 3400
rect 4250 2800 4310 3400
rect 4590 2800 4650 3400
rect 5050 2800 5110 3400
rect 5390 2800 5450 3400
rect 5850 2800 5910 3400
rect 6190 2800 6250 3400
rect 6650 2800 6710 3400
rect 6990 2800 7050 3400
rect 7450 2800 7510 3400
rect 7790 2800 7850 3400
rect 8250 2800 8310 3400
rect 8590 2800 8650 3400
rect 9050 2800 9110 3400
rect 9390 2800 9450 3400
rect 9850 2800 9910 3400
rect 10190 2800 10250 3400
rect 10650 2800 10710 3400
rect 10990 2800 11050 3400
rect 11450 2800 11510 3400
rect 11790 2800 11850 3400
rect 12250 2800 12310 3400
rect 12590 2800 12650 3400
rect 250 2000 310 2600
rect 590 2000 650 2600
rect 1050 2000 1110 2600
rect 1390 2000 1450 2600
rect 1850 2000 1910 2600
rect 2190 2000 2250 2600
rect 2650 2000 2710 2600
rect 2990 2000 3050 2600
rect 3450 2000 3510 2600
rect 3790 2000 3850 2600
rect 4250 2000 4310 2600
rect 4590 2000 4650 2600
rect 5050 2000 5110 2600
rect 5390 2000 5450 2600
rect 5850 2000 5910 2600
rect 6190 2000 6250 2600
rect 6650 2000 6710 2600
rect 6990 2000 7050 2600
rect 7450 2000 7510 2600
rect 7790 2000 7850 2600
rect 8250 2000 8310 2600
rect 8590 2000 8650 2600
rect 9050 2000 9110 2600
rect 9390 2000 9450 2600
rect 9850 2000 9910 2600
rect 10190 2000 10250 2600
rect 10650 2000 10710 2600
rect 10990 2000 11050 2600
rect 11450 2000 11510 2600
rect 11790 2000 11850 2600
rect 12250 2000 12310 2600
rect 12590 2000 12650 2600
rect 250 1200 310 1800
rect 590 1200 650 1800
rect 1050 1200 1110 1800
rect 1390 1200 1450 1800
rect 1850 1200 1910 1800
rect 2190 1200 2250 1800
rect 2650 1200 2710 1800
rect 2990 1200 3050 1800
rect 3450 1200 3510 1800
rect 3790 1200 3850 1800
rect 4250 1200 4310 1800
rect 4590 1200 4650 1800
rect 5050 1200 5110 1800
rect 5390 1200 5450 1800
rect 5850 1200 5910 1800
rect 6190 1200 6250 1800
rect 6650 1200 6710 1800
rect 6990 1200 7050 1800
rect 7450 1200 7510 1800
rect 7790 1200 7850 1800
rect 8250 1200 8310 1800
rect 8590 1200 8650 1800
rect 9050 1200 9110 1800
rect 9390 1200 9450 1800
rect 9850 1200 9910 1800
rect 10190 1200 10250 1800
rect 10650 1200 10710 1800
rect 10990 1200 11050 1800
rect 11450 1200 11510 1800
rect 11790 1200 11850 1800
rect 12250 1200 12310 1800
rect 12590 1200 12650 1800
rect 250 400 310 1000
rect 590 400 650 1000
rect 1050 400 1110 1000
rect 1390 400 1450 1000
rect 1850 400 1910 1000
rect 2190 400 2250 1000
rect 2650 400 2710 1000
rect 2990 400 3050 1000
rect 3450 400 3510 1000
rect 3790 400 3850 1000
rect 4250 400 4310 1000
rect 4590 400 4650 1000
rect 5050 400 5110 1000
rect 5390 400 5450 1000
rect 5850 400 5910 1000
rect 6190 400 6250 1000
rect 6650 400 6710 1000
rect 6990 400 7050 1000
rect 7450 400 7510 1000
rect 7790 400 7850 1000
rect 8250 400 8310 1000
rect 8590 400 8650 1000
rect 9050 400 9110 1000
rect 9390 400 9450 1000
rect 9850 400 9910 1000
rect 10190 400 10250 1000
rect 10650 400 10710 1000
rect 10990 400 11050 1000
rect 11450 400 11510 1000
rect 11790 400 11850 1000
rect 12250 400 12310 1000
rect 12590 400 12650 1000
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
array 0 15 800 0 7 800
timestamp 1667663783
transform 1 0 325 0 1 300
box -325 -300 325 300
<< end >>
