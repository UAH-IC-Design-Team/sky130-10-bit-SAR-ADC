magic
tech sky130A
magscale 1 2
timestamp 1666486738
<< error_p >>
rect -29 2227 29 2233
rect -29 2193 -17 2227
rect -29 2187 29 2193
rect -29 1769 29 1775
rect -29 1735 -17 1769
rect -29 1729 29 1735
rect -29 1661 29 1667
rect -29 1627 -17 1661
rect -29 1621 29 1627
rect -29 1203 29 1209
rect -29 1169 -17 1203
rect -29 1163 29 1169
rect -29 1095 29 1101
rect -29 1061 -17 1095
rect -29 1055 29 1061
rect -29 637 29 643
rect -29 603 -17 637
rect -29 597 29 603
rect -29 529 29 535
rect -29 495 -17 529
rect -29 489 29 495
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -495 29 -489
rect -29 -529 -17 -495
rect -29 -535 29 -529
rect -29 -603 29 -597
rect -29 -637 -17 -603
rect -29 -643 29 -637
rect -29 -1061 29 -1055
rect -29 -1095 -17 -1061
rect -29 -1101 29 -1095
rect -29 -1169 29 -1163
rect -29 -1203 -17 -1169
rect -29 -1209 29 -1203
rect -29 -1627 29 -1621
rect -29 -1661 -17 -1627
rect -29 -1667 29 -1661
rect -29 -1735 29 -1729
rect -29 -1769 -17 -1735
rect -29 -1775 29 -1769
rect -29 -2193 29 -2187
rect -29 -2227 -17 -2193
rect -29 -2233 29 -2227
<< nwell >>
rect -211 -2365 211 2365
<< pmos >>
rect -15 1816 15 2146
rect -15 1250 15 1580
rect -15 684 15 1014
rect -15 118 15 448
rect -15 -448 15 -118
rect -15 -1014 15 -684
rect -15 -1580 15 -1250
rect -15 -2146 15 -1816
<< pdiff >>
rect -73 2134 -15 2146
rect -73 1828 -61 2134
rect -27 1828 -15 2134
rect -73 1816 -15 1828
rect 15 2134 73 2146
rect 15 1828 27 2134
rect 61 1828 73 2134
rect 15 1816 73 1828
rect -73 1568 -15 1580
rect -73 1262 -61 1568
rect -27 1262 -15 1568
rect -73 1250 -15 1262
rect 15 1568 73 1580
rect 15 1262 27 1568
rect 61 1262 73 1568
rect 15 1250 73 1262
rect -73 1002 -15 1014
rect -73 696 -61 1002
rect -27 696 -15 1002
rect -73 684 -15 696
rect 15 1002 73 1014
rect 15 696 27 1002
rect 61 696 73 1002
rect 15 684 73 696
rect -73 436 -15 448
rect -73 130 -61 436
rect -27 130 -15 436
rect -73 118 -15 130
rect 15 436 73 448
rect 15 130 27 436
rect 61 130 73 436
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -436 -61 -130
rect -27 -436 -15 -130
rect -73 -448 -15 -436
rect 15 -130 73 -118
rect 15 -436 27 -130
rect 61 -436 73 -130
rect 15 -448 73 -436
rect -73 -696 -15 -684
rect -73 -1002 -61 -696
rect -27 -1002 -15 -696
rect -73 -1014 -15 -1002
rect 15 -696 73 -684
rect 15 -1002 27 -696
rect 61 -1002 73 -696
rect 15 -1014 73 -1002
rect -73 -1262 -15 -1250
rect -73 -1568 -61 -1262
rect -27 -1568 -15 -1262
rect -73 -1580 -15 -1568
rect 15 -1262 73 -1250
rect 15 -1568 27 -1262
rect 61 -1568 73 -1262
rect 15 -1580 73 -1568
rect -73 -1828 -15 -1816
rect -73 -2134 -61 -1828
rect -27 -2134 -15 -1828
rect -73 -2146 -15 -2134
rect 15 -1828 73 -1816
rect 15 -2134 27 -1828
rect 61 -2134 73 -1828
rect 15 -2146 73 -2134
<< pdiffc >>
rect -61 1828 -27 2134
rect 27 1828 61 2134
rect -61 1262 -27 1568
rect 27 1262 61 1568
rect -61 696 -27 1002
rect 27 696 61 1002
rect -61 130 -27 436
rect 27 130 61 436
rect -61 -436 -27 -130
rect 27 -436 61 -130
rect -61 -1002 -27 -696
rect 27 -1002 61 -696
rect -61 -1568 -27 -1262
rect 27 -1568 61 -1262
rect -61 -2134 -27 -1828
rect 27 -2134 61 -1828
<< nsubdiff >>
rect -175 2295 -79 2329
rect 79 2295 175 2329
rect -175 2233 -141 2295
rect 141 2233 175 2295
rect -175 -2295 -141 -2233
rect 141 -2295 175 -2233
rect -175 -2329 -79 -2295
rect 79 -2329 175 -2295
<< nsubdiffcont >>
rect -79 2295 79 2329
rect -175 -2233 -141 2233
rect 141 -2233 175 2233
rect -79 -2329 79 -2295
<< poly >>
rect -33 2227 33 2243
rect -33 2193 -17 2227
rect 17 2193 33 2227
rect -33 2177 33 2193
rect -15 2146 15 2177
rect -15 1785 15 1816
rect -33 1769 33 1785
rect -33 1735 -17 1769
rect 17 1735 33 1769
rect -33 1719 33 1735
rect -33 1661 33 1677
rect -33 1627 -17 1661
rect 17 1627 33 1661
rect -33 1611 33 1627
rect -15 1580 15 1611
rect -15 1219 15 1250
rect -33 1203 33 1219
rect -33 1169 -17 1203
rect 17 1169 33 1203
rect -33 1153 33 1169
rect -33 1095 33 1111
rect -33 1061 -17 1095
rect 17 1061 33 1095
rect -33 1045 33 1061
rect -15 1014 15 1045
rect -15 653 15 684
rect -33 637 33 653
rect -33 603 -17 637
rect 17 603 33 637
rect -33 587 33 603
rect -33 529 33 545
rect -33 495 -17 529
rect 17 495 33 529
rect -33 479 33 495
rect -15 448 15 479
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -479 15 -448
rect -33 -495 33 -479
rect -33 -529 -17 -495
rect 17 -529 33 -495
rect -33 -545 33 -529
rect -33 -603 33 -587
rect -33 -637 -17 -603
rect 17 -637 33 -603
rect -33 -653 33 -637
rect -15 -684 15 -653
rect -15 -1045 15 -1014
rect -33 -1061 33 -1045
rect -33 -1095 -17 -1061
rect 17 -1095 33 -1061
rect -33 -1111 33 -1095
rect -33 -1169 33 -1153
rect -33 -1203 -17 -1169
rect 17 -1203 33 -1169
rect -33 -1219 33 -1203
rect -15 -1250 15 -1219
rect -15 -1611 15 -1580
rect -33 -1627 33 -1611
rect -33 -1661 -17 -1627
rect 17 -1661 33 -1627
rect -33 -1677 33 -1661
rect -33 -1735 33 -1719
rect -33 -1769 -17 -1735
rect 17 -1769 33 -1735
rect -33 -1785 33 -1769
rect -15 -1816 15 -1785
rect -15 -2177 15 -2146
rect -33 -2193 33 -2177
rect -33 -2227 -17 -2193
rect 17 -2227 33 -2193
rect -33 -2243 33 -2227
<< polycont >>
rect -17 2193 17 2227
rect -17 1735 17 1769
rect -17 1627 17 1661
rect -17 1169 17 1203
rect -17 1061 17 1095
rect -17 603 17 637
rect -17 495 17 529
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -529 17 -495
rect -17 -637 17 -603
rect -17 -1095 17 -1061
rect -17 -1203 17 -1169
rect -17 -1661 17 -1627
rect -17 -1769 17 -1735
rect -17 -2227 17 -2193
<< locali >>
rect -175 2295 -79 2329
rect 79 2295 175 2329
rect -175 2233 -141 2295
rect 141 2233 175 2295
rect -33 2193 -17 2227
rect 17 2193 33 2227
rect -61 2134 -27 2150
rect -61 1812 -27 1828
rect 27 2134 61 2150
rect 27 1812 61 1828
rect -33 1735 -17 1769
rect 17 1735 33 1769
rect -33 1627 -17 1661
rect 17 1627 33 1661
rect -61 1568 -27 1584
rect -61 1246 -27 1262
rect 27 1568 61 1584
rect 27 1246 61 1262
rect -33 1169 -17 1203
rect 17 1169 33 1203
rect -33 1061 -17 1095
rect 17 1061 33 1095
rect -61 1002 -27 1018
rect -61 680 -27 696
rect 27 1002 61 1018
rect 27 680 61 696
rect -33 603 -17 637
rect 17 603 33 637
rect -33 495 -17 529
rect 17 495 33 529
rect -61 436 -27 452
rect -61 114 -27 130
rect 27 436 61 452
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -452 -27 -436
rect 27 -130 61 -114
rect 27 -452 61 -436
rect -33 -529 -17 -495
rect 17 -529 33 -495
rect -33 -637 -17 -603
rect 17 -637 33 -603
rect -61 -696 -27 -680
rect -61 -1018 -27 -1002
rect 27 -696 61 -680
rect 27 -1018 61 -1002
rect -33 -1095 -17 -1061
rect 17 -1095 33 -1061
rect -33 -1203 -17 -1169
rect 17 -1203 33 -1169
rect -61 -1262 -27 -1246
rect -61 -1584 -27 -1568
rect 27 -1262 61 -1246
rect 27 -1584 61 -1568
rect -33 -1661 -17 -1627
rect 17 -1661 33 -1627
rect -33 -1769 -17 -1735
rect 17 -1769 33 -1735
rect -61 -1828 -27 -1812
rect -61 -2150 -27 -2134
rect 27 -1828 61 -1812
rect 27 -2150 61 -2134
rect -33 -2227 -17 -2193
rect 17 -2227 33 -2193
rect -175 -2295 -141 -2233
rect 141 -2295 175 -2233
rect -175 -2329 -79 -2295
rect 79 -2329 175 -2295
<< viali >>
rect -17 2193 17 2227
rect -61 1828 -27 2134
rect 27 1828 61 2134
rect -17 1735 17 1769
rect -17 1627 17 1661
rect -61 1262 -27 1568
rect 27 1262 61 1568
rect -17 1169 17 1203
rect -17 1061 17 1095
rect -61 696 -27 1002
rect 27 696 61 1002
rect -17 603 17 637
rect -17 495 17 529
rect -61 130 -27 436
rect 27 130 61 436
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -436 -27 -130
rect 27 -436 61 -130
rect -17 -529 17 -495
rect -17 -637 17 -603
rect -61 -1002 -27 -696
rect 27 -1002 61 -696
rect -17 -1095 17 -1061
rect -17 -1203 17 -1169
rect -61 -1568 -27 -1262
rect 27 -1568 61 -1262
rect -17 -1661 17 -1627
rect -17 -1769 17 -1735
rect -61 -2134 -27 -1828
rect 27 -2134 61 -1828
rect -17 -2227 17 -2193
<< metal1 >>
rect -29 2227 29 2233
rect -29 2193 -17 2227
rect 17 2193 29 2227
rect -29 2187 29 2193
rect -67 2134 -21 2146
rect -67 1828 -61 2134
rect -27 1828 -21 2134
rect -67 1816 -21 1828
rect 21 2134 67 2146
rect 21 1828 27 2134
rect 61 1828 67 2134
rect 21 1816 67 1828
rect -29 1769 29 1775
rect -29 1735 -17 1769
rect 17 1735 29 1769
rect -29 1729 29 1735
rect -29 1661 29 1667
rect -29 1627 -17 1661
rect 17 1627 29 1661
rect -29 1621 29 1627
rect -67 1568 -21 1580
rect -67 1262 -61 1568
rect -27 1262 -21 1568
rect -67 1250 -21 1262
rect 21 1568 67 1580
rect 21 1262 27 1568
rect 61 1262 67 1568
rect 21 1250 67 1262
rect -29 1203 29 1209
rect -29 1169 -17 1203
rect 17 1169 29 1203
rect -29 1163 29 1169
rect -29 1095 29 1101
rect -29 1061 -17 1095
rect 17 1061 29 1095
rect -29 1055 29 1061
rect -67 1002 -21 1014
rect -67 696 -61 1002
rect -27 696 -21 1002
rect -67 684 -21 696
rect 21 1002 67 1014
rect 21 696 27 1002
rect 61 696 67 1002
rect 21 684 67 696
rect -29 637 29 643
rect -29 603 -17 637
rect 17 603 29 637
rect -29 597 29 603
rect -29 529 29 535
rect -29 495 -17 529
rect 17 495 29 529
rect -29 489 29 495
rect -67 436 -21 448
rect -67 130 -61 436
rect -27 130 -21 436
rect -67 118 -21 130
rect 21 436 67 448
rect 21 130 27 436
rect 61 130 67 436
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -436 -61 -130
rect -27 -436 -21 -130
rect -67 -448 -21 -436
rect 21 -130 67 -118
rect 21 -436 27 -130
rect 61 -436 67 -130
rect 21 -448 67 -436
rect -29 -495 29 -489
rect -29 -529 -17 -495
rect 17 -529 29 -495
rect -29 -535 29 -529
rect -29 -603 29 -597
rect -29 -637 -17 -603
rect 17 -637 29 -603
rect -29 -643 29 -637
rect -67 -696 -21 -684
rect -67 -1002 -61 -696
rect -27 -1002 -21 -696
rect -67 -1014 -21 -1002
rect 21 -696 67 -684
rect 21 -1002 27 -696
rect 61 -1002 67 -696
rect 21 -1014 67 -1002
rect -29 -1061 29 -1055
rect -29 -1095 -17 -1061
rect 17 -1095 29 -1061
rect -29 -1101 29 -1095
rect -29 -1169 29 -1163
rect -29 -1203 -17 -1169
rect 17 -1203 29 -1169
rect -29 -1209 29 -1203
rect -67 -1262 -21 -1250
rect -67 -1568 -61 -1262
rect -27 -1568 -21 -1262
rect -67 -1580 -21 -1568
rect 21 -1262 67 -1250
rect 21 -1568 27 -1262
rect 61 -1568 67 -1262
rect 21 -1580 67 -1568
rect -29 -1627 29 -1621
rect -29 -1661 -17 -1627
rect 17 -1661 29 -1627
rect -29 -1667 29 -1661
rect -29 -1735 29 -1729
rect -29 -1769 -17 -1735
rect 17 -1769 29 -1735
rect -29 -1775 29 -1769
rect -67 -1828 -21 -1816
rect -67 -2134 -61 -1828
rect -27 -2134 -21 -1828
rect -67 -2146 -21 -2134
rect 21 -1828 67 -1816
rect 21 -2134 27 -1828
rect 61 -2134 67 -1828
rect 21 -2146 67 -2134
rect -29 -2193 29 -2187
rect -29 -2227 -17 -2193
rect 17 -2227 29 -2193
rect -29 -2233 29 -2227
<< properties >>
string FIXED_BBOX -158 -2312 158 2312
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
