magic
tech sky130A
magscale 1 2
timestamp 1666918578
<< error_p >>
rect -77 242 -19 248
rect 115 242 173 248
rect -77 208 -65 242
rect 115 208 127 242
rect -77 202 -19 208
rect 115 202 173 208
rect -173 -208 -115 -202
rect 19 -208 77 -202
rect -173 -242 -161 -208
rect 19 -242 31 -208
rect -173 -248 -115 -242
rect 19 -248 77 -242
<< nwell >>
rect -161 223 257 261
rect -257 -223 257 223
rect -257 -261 161 -223
<< pmos >>
rect -159 -161 -129 161
rect -63 -161 -33 161
rect 33 -161 63 161
rect 129 -161 159 161
<< pdiff >>
rect -221 149 -159 161
rect -221 -149 -209 149
rect -175 -149 -159 149
rect -221 -161 -159 -149
rect -129 149 -63 161
rect -129 -149 -113 149
rect -79 -149 -63 149
rect -129 -161 -63 -149
rect -33 149 33 161
rect -33 -149 -17 149
rect 17 -149 33 149
rect -33 -161 33 -149
rect 63 149 129 161
rect 63 -149 79 149
rect 113 -149 129 149
rect 63 -161 129 -149
rect 159 149 221 161
rect 159 -149 175 149
rect 209 -149 221 149
rect 159 -161 221 -149
<< pdiffc >>
rect -209 -149 -175 149
rect -113 -149 -79 149
rect -17 -149 17 149
rect 79 -149 113 149
rect 175 -149 209 149
<< poly >>
rect -81 242 -15 258
rect -81 208 -65 242
rect -31 208 -15 242
rect -81 192 -15 208
rect 111 242 177 258
rect 111 208 127 242
rect 161 208 177 242
rect 111 192 177 208
rect -159 161 -129 187
rect -63 161 -33 192
rect 33 161 63 187
rect 129 161 159 192
rect -159 -192 -129 -161
rect -63 -187 -33 -161
rect 33 -192 63 -161
rect 129 -187 159 -161
rect -177 -208 -111 -192
rect -177 -242 -161 -208
rect -127 -242 -111 -208
rect -177 -258 -111 -242
rect 15 -208 81 -192
rect 15 -242 31 -208
rect 65 -242 81 -208
rect 15 -258 81 -242
<< polycont >>
rect -65 208 -31 242
rect 127 208 161 242
rect -161 -242 -127 -208
rect 31 -242 65 -208
<< locali >>
rect -81 208 -65 242
rect -31 208 -15 242
rect 111 208 127 242
rect 161 208 177 242
rect -209 149 -175 165
rect -209 -165 -175 -149
rect -113 149 -79 165
rect -113 -165 -79 -149
rect -17 149 17 165
rect -17 -165 17 -149
rect 79 149 113 165
rect 79 -165 113 -149
rect 175 149 209 165
rect 175 -165 209 -149
rect -177 -242 -161 -208
rect -127 -242 -111 -208
rect 15 -242 31 -208
rect 65 -242 81 -208
<< viali >>
rect -65 208 -31 242
rect 127 208 161 242
rect -209 -149 -175 149
rect -113 -149 -79 149
rect -17 -149 17 149
rect 79 -149 113 149
rect 175 -149 209 149
rect -161 -242 -127 -208
rect 31 -242 65 -208
<< metal1 >>
rect -77 242 -19 248
rect -77 208 -65 242
rect -31 208 -19 242
rect -77 202 -19 208
rect 115 242 173 248
rect 115 208 127 242
rect 161 208 173 242
rect 115 202 173 208
rect -215 149 -169 161
rect -215 -149 -209 149
rect -175 -149 -169 149
rect -215 -161 -169 -149
rect -119 149 -73 161
rect -119 -149 -113 149
rect -79 -149 -73 149
rect -119 -161 -73 -149
rect -23 149 23 161
rect -23 -149 -17 149
rect 17 -149 23 149
rect -23 -161 23 -149
rect 73 149 119 161
rect 73 -149 79 149
rect 113 -149 119 149
rect 73 -161 119 -149
rect 169 149 215 161
rect 169 -149 175 149
rect 209 -149 215 149
rect 169 -161 215 -149
rect -173 -208 -115 -202
rect -173 -242 -161 -208
rect -127 -242 -115 -208
rect -173 -248 -115 -242
rect 19 -208 77 -202
rect 19 -242 31 -208
rect 65 -242 77 -208
rect 19 -248 77 -242
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
