magic
tech sky130A
magscale 1 2
timestamp 1666292354
<< metal3 >>
rect -892 2117 -120 2145
rect -892 -2117 -204 2117
rect -140 -2117 -120 2117
rect -892 -2145 -120 -2117
rect 120 2117 892 2145
rect 120 -2117 808 2117
rect 872 -2117 892 2117
rect 120 -2145 892 -2117
<< via3 >>
rect -204 -2117 -140 2117
rect 808 -2117 872 2117
<< mimcap >>
rect -852 2065 -452 2105
rect -852 -2065 -812 2065
rect -492 -2065 -452 2065
rect -852 -2105 -452 -2065
rect 160 2065 560 2105
rect 160 -2065 200 2065
rect 520 -2065 560 2065
rect 160 -2105 560 -2065
<< mimcapcontact >>
rect -812 -2065 -492 2065
rect 200 -2065 520 2065
<< metal4 >>
rect -220 2117 -124 2133
rect -813 2065 -491 2066
rect -813 -2065 -812 2065
rect -492 -2065 -491 2065
rect -813 -2066 -491 -2065
rect -220 -2117 -204 2117
rect -140 -2117 -124 2117
rect 792 2117 888 2133
rect 199 2065 521 2066
rect 199 -2065 200 2065
rect 520 -2065 521 2065
rect 199 -2066 521 -2065
rect -220 -2133 -124 -2117
rect 792 -2117 808 2117
rect 872 -2117 888 2117
rect 792 -2133 888 -2117
<< properties >>
string FIXED_BBOX 120 -2145 600 2145
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 21.052 val 92.967 carea 2.00 cperi 0.19 nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
