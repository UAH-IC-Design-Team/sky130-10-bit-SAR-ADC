** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/tests/demux2/demux2_test.sch
**.subckt demux2_test
V3 VDD GND 1.8V
V4 VSS GND 0
x1 select out_0 v_in out_1 VDD VSS demux2
V1 select GND PULSE 0 1.8V 0 1ns 1ns 10us 20us
V2 v_in GND PULSE 0 1.8V 0 1ns 1ns 7us 15us
**** begin user architecture code
* .lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* .include /foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


.options acct list
.temp 25
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
.control
tran 0.1u 100u
plot select v_in+2 out_0+4 out_1+6
write dmux2_test_with_xspice.raw
.endc



* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sch

* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sch
.subckt demux2 a_S a_OUT_0 a_IN a_OUT_1 a_VDD a_VSS
*.PININFO S:I OUT_0:O IN:I OUT_1:O VDD:B VSS:B
A1 [net1 IN] OUT_0 d_lut_sky130_fd_sc_hd__and2_0
A2 [S IN] OUT_1 d_lut_sky130_fd_sc_hd__and2_0
A3 [S] net1 d_lut_sky130_fd_sc_hd__inv_1
**** begin user architecture code
**** end user architecture code

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_S] [S] todig_1v8
AD2A1 [OUT_0] [a_OUT_0] toana_1v8
AA2D2 [a_IN] [IN] todig_1v8
AD2A2 [OUT_1] [a_OUT_1] toana_1v8
AA2D3 [a_VDD] [VDD] todig_1v8
AA2D4 [a_VSS] [VSS] todig_1v8

.ends

* sky130_fd_sc_hd__and2_0 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_0 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__inv_1 (!A)
.model d_lut_sky130_fd_sc_hd__inv_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10")

.GLOBAL GND
.end
