magic
tech sky130A
magscale 1 2
timestamp 1666649035
<< error_p >>
rect -29 242 29 248
rect -29 208 -17 242
rect -29 202 29 208
rect -29 -208 29 -202
rect -29 -242 -17 -208
rect -29 -248 29 -242
<< nwell >>
rect -211 -380 211 380
<< pmos >>
rect -15 -161 15 161
<< pdiff >>
rect -73 149 -15 161
rect -73 -149 -61 149
rect -27 -149 -15 149
rect -73 -161 -15 -149
rect 15 149 73 161
rect 15 -149 27 149
rect 61 -149 73 149
rect 15 -161 73 -149
<< pdiffc >>
rect -61 -149 -27 149
rect 27 -149 61 149
<< nsubdiff >>
rect -175 310 -79 344
rect 79 310 175 344
rect -175 248 -141 310
rect 141 248 175 310
rect -175 -310 -141 -248
rect 141 -310 175 -248
rect -175 -344 -79 -310
rect 79 -344 175 -310
<< nsubdiffcont >>
rect -79 310 79 344
rect -175 -248 -141 248
rect 141 -248 175 248
rect -79 -344 79 -310
<< poly >>
rect -33 242 33 258
rect -33 208 -17 242
rect 17 208 33 242
rect -33 192 33 208
rect -15 161 15 192
rect -15 -192 15 -161
rect -33 -208 33 -192
rect -33 -242 -17 -208
rect 17 -242 33 -208
rect -33 -258 33 -242
<< polycont >>
rect -17 208 17 242
rect -17 -242 17 -208
<< locali >>
rect -175 310 -79 344
rect 79 310 175 344
rect -175 248 -141 310
rect 141 248 175 310
rect -33 208 -17 242
rect 17 208 33 242
rect -61 149 -27 165
rect -61 -165 -27 -149
rect 27 149 61 165
rect 27 -165 61 -149
rect -33 -242 -17 -208
rect 17 -242 33 -208
rect -175 -310 -141 -248
rect 141 -310 175 -248
rect -175 -344 -79 -310
rect 79 -344 175 -310
<< viali >>
rect -17 208 17 242
rect -61 -149 -27 149
rect 27 -149 61 149
rect -17 -242 17 -208
<< metal1 >>
rect -29 242 29 248
rect -29 208 -17 242
rect 17 208 29 242
rect -29 202 29 208
rect -67 149 -21 161
rect -67 -149 -61 149
rect -27 -149 -21 149
rect -67 -161 -21 -149
rect 21 149 67 161
rect 21 -149 27 149
rect 61 -149 67 149
rect 21 -161 67 -149
rect -29 -208 29 -202
rect -29 -242 -17 -208
rect 17 -242 29 -208
rect -29 -248 29 -242
<< properties >>
string FIXED_BBOX -158 -327 158 327
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.605 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
