magic
tech sky130A
magscale 1 2
timestamp 1667500205
<< error_p >>
rect -269 222 -207 1000
rect -177 222 -111 1000
rect -81 222 -15 1000
rect 15 222 81 1000
rect 111 222 177 1000
rect 207 222 269 1000
<< nmos >>
rect -207 -1000 -177 1000
rect -111 -1000 -81 1000
rect -15 -1000 15 1000
rect 81 -1000 111 1000
rect 177 -1000 207 1000
<< ndiff >>
rect -269 988 -207 1000
rect -269 -988 -257 988
rect -223 -988 -207 988
rect -269 -1000 -207 -988
rect -177 988 -111 1000
rect -177 -988 -161 988
rect -127 -988 -111 988
rect -177 -1000 -111 -988
rect -81 988 -15 1000
rect -81 -988 -65 988
rect -31 -988 -15 988
rect -81 -1000 -15 -988
rect 15 988 81 1000
rect 15 -988 31 988
rect 65 -988 81 988
rect 15 -1000 81 -988
rect 111 988 177 1000
rect 111 -988 127 988
rect 161 -988 177 988
rect 111 -1000 177 -988
rect 207 988 269 1000
rect 207 -988 223 988
rect 257 -988 269 988
rect 207 -1000 269 -988
<< ndiffc >>
rect -257 -988 -223 988
rect -161 -988 -127 988
rect -65 -988 -31 988
rect 31 -988 65 988
rect 127 -988 161 988
rect 223 -988 257 988
<< poly >>
rect -207 1000 -177 1028
rect -111 1000 -81 1028
rect -15 1000 15 1028
rect 81 1000 111 1028
rect 177 1000 207 1028
rect -207 -1022 -177 -1000
rect -111 -1022 -81 -1000
rect -15 -1022 15 -1000
rect 81 -1022 111 -1000
rect 177 -1022 207 -1000
rect -225 -1038 231 -1022
rect -225 -1072 -209 -1038
rect -175 -1072 -114 -1038
rect -80 -1072 -17 -1038
rect 17 -1072 76 -1038
rect 110 -1072 175 -1038
rect 209 -1072 231 -1038
rect -225 -1088 231 -1072
<< polycont >>
rect -209 -1072 -175 -1038
rect -114 -1072 -80 -1038
rect -17 -1072 17 -1038
rect 76 -1072 110 -1038
rect 175 -1072 209 -1038
<< locali >>
rect -257 988 -223 1004
rect -257 -1004 -223 -988
rect -161 988 -127 1004
rect -161 -1004 -127 -988
rect -65 988 -31 1004
rect -65 -1004 -31 -988
rect 31 988 65 1004
rect 31 -1004 65 -988
rect 127 988 161 1004
rect 127 -1004 161 -988
rect 223 988 257 1004
rect 223 -1004 257 -988
rect -225 -1072 -209 -1038
rect -175 -1072 -114 -1038
rect -80 -1072 -17 -1038
rect 17 -1072 76 -1038
rect 110 -1072 175 -1038
rect 209 -1072 231 -1038
<< viali >>
rect -257 -971 -223 -181
rect -161 181 -127 971
rect -65 -971 -31 -181
rect 31 181 65 971
rect 127 -971 161 -181
rect 223 181 257 971
rect -209 -1072 -175 -1038
rect -114 -1072 -80 -1038
rect -17 -1072 17 -1038
rect 76 -1072 110 -1038
rect 175 -1072 209 -1038
<< metal1 >>
rect -167 971 -121 983
rect -167 181 -161 971
rect -127 181 -121 971
rect -167 169 -121 181
rect 25 971 71 983
rect 25 181 31 971
rect 65 181 71 971
rect 25 169 71 181
rect 217 971 263 983
rect 217 181 223 971
rect 257 181 263 971
rect 217 169 263 181
rect -263 -181 -217 -169
rect -263 -971 -257 -181
rect -223 -971 -217 -181
rect -263 -983 -217 -971
rect -71 -181 -25 -169
rect -71 -971 -65 -181
rect -31 -971 -25 -181
rect -71 -983 -25 -971
rect 121 -181 167 -169
rect 121 -971 127 -181
rect 161 -971 167 -181
rect 121 -983 167 -971
rect -225 -1038 231 -1032
rect -225 -1072 -209 -1038
rect -175 -1072 -114 -1038
rect -80 -1072 -17 -1038
rect 17 -1072 76 -1038
rect 110 -1072 175 -1038
rect 209 -1072 231 -1038
rect -225 -1078 231 -1072
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
