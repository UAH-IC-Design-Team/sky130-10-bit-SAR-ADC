* XSpice netlist created from SPICE and liberty sources by spi2xspice.py
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/tests/demux2/demux2_test.sch
**.subckt demux2_test
**** begin user architecture code
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
**** end user architecture code
**.ends
* expanding   symbol:  src/demux2/demux2.sym # of pins=6
** sym_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sym
** sch_path: /foss/designs/sky130-10-bit-SAR-ADC/xschem/src/demux2/demux2.sch
.subckt demux2 a_S a_VDD a_VSS a_OUT_0 a_IN a_OUT_1
*.ipin S
*.opin OUT_0
*.ipin IN
*.opin OUT_1
*.iopin VDD
*.iopin VSS
A1 [net1 IN] OUT_0 d_lut_sky130_fd_sc_hd__and2_0
A2 [S IN] OUT_1 d_lut_sky130_fd_sc_hd__and2_0
A3 [S] net1 d_lut_sky130_fd_sc_hd__inv_1

.model todig_1v8 adc_bridge(in_high=1.2 in_low=0.6 rise_delay=10n fall_delay=10n)
.model toana_1v8 dac_bridge(out_high=1.8 out_low=0)

.model ddflop d_dff(ic=0 rise_delay=1n fall_delay=1n)
.model dzero d_pulldown(load=1p)
.model done d_pullup(load=1p)

AA2D1 [a_S] [S] todig_1v8
AA2D2 [a_VDD] [VDD] todig_1v8
AA2D3 [a_VSS] [VSS] todig_1v8
AD2A1 [OUT_0] [a_OUT_0] toana_1v8
AA2D4 [a_IN] [IN] todig_1v8
AD2A2 [OUT_1] [a_OUT_1] toana_1v8

.ends

.GLOBAL GND

* sky130_fd_sc_hd__and2_0 (A&B)
.model d_lut_sky130_fd_sc_hd__and2_0 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "0001")
* sky130_fd_sc_hd__inv_1 (!A)
.model d_lut_sky130_fd_sc_hd__inv_1 d_lut (rise_delay=1n fall_delay=1n input_load=1p
+ table_values "10")
.end
