magic
tech sky130A
magscale 1 2
timestamp 1666552007
<< error_p >>
rect -29 4491 29 4497
rect -29 4457 -17 4491
rect -29 4451 29 4457
rect -109 3980 109 4198
rect -29 3925 29 3931
rect -29 3891 -17 3925
rect -29 3885 29 3891
rect -109 3414 109 3632
rect -29 3359 29 3365
rect -29 3325 -17 3359
rect -29 3319 29 3325
rect -109 2848 109 3066
rect -29 2793 29 2799
rect -29 2759 -17 2793
rect -29 2753 29 2759
rect -109 2282 109 2500
rect -29 2227 29 2233
rect -29 2193 -17 2227
rect -29 2187 29 2193
rect -109 1716 109 1934
rect -29 1661 29 1667
rect -29 1627 -17 1661
rect -29 1621 29 1627
rect -109 1150 109 1368
rect -29 1095 29 1101
rect -29 1061 -17 1095
rect -29 1055 29 1061
rect -109 584 109 802
rect -29 529 29 535
rect -29 495 -17 529
rect -29 489 29 495
rect -109 18 109 236
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -109 -548 109 -330
rect -29 -603 29 -597
rect -29 -637 -17 -603
rect -29 -643 29 -637
rect -109 -1114 109 -896
rect -29 -1169 29 -1163
rect -29 -1203 -17 -1169
rect -29 -1209 29 -1203
rect -109 -1680 109 -1462
rect -29 -1735 29 -1729
rect -29 -1769 -17 -1735
rect -29 -1775 29 -1769
rect -109 -2246 109 -2028
rect -29 -2301 29 -2295
rect -29 -2335 -17 -2301
rect -29 -2341 29 -2335
rect -109 -2812 109 -2594
rect -29 -2867 29 -2861
rect -29 -2901 -17 -2867
rect -29 -2907 29 -2901
rect -109 -3378 109 -3160
rect -29 -3433 29 -3427
rect -29 -3467 -17 -3433
rect -29 -3473 29 -3467
rect -109 -3944 109 -3726
rect -29 -3999 29 -3993
rect -29 -4033 -17 -3999
rect -29 -4039 29 -4033
rect -29 -4457 29 -4451
rect -29 -4491 -17 -4457
rect -29 -4497 29 -4491
<< nwell >>
rect -109 3980 109 4510
rect -109 3414 109 3944
rect -109 2848 109 3378
rect -109 2282 109 2812
rect -109 1716 109 2246
rect -109 1150 109 1680
rect -109 584 109 1114
rect -109 18 109 548
rect -109 -548 109 -18
rect -109 -1114 109 -584
rect -109 -1680 109 -1150
rect -109 -2246 109 -1716
rect -109 -2812 109 -2282
rect -109 -3378 109 -2848
rect -109 -3944 109 -3414
rect -109 -4510 109 -3980
<< pmos >>
rect -15 4080 15 4410
rect -15 3514 15 3844
rect -15 2948 15 3278
rect -15 2382 15 2712
rect -15 1816 15 2146
rect -15 1250 15 1580
rect -15 684 15 1014
rect -15 118 15 448
rect -15 -448 15 -118
rect -15 -1014 15 -684
rect -15 -1580 15 -1250
rect -15 -2146 15 -1816
rect -15 -2712 15 -2382
rect -15 -3278 15 -2948
rect -15 -3844 15 -3514
rect -15 -4410 15 -4080
<< pdiff >>
rect -73 4398 -15 4410
rect -73 4092 -61 4398
rect -27 4092 -15 4398
rect -73 4080 -15 4092
rect 15 4398 73 4410
rect 15 4092 27 4398
rect 61 4092 73 4398
rect 15 4080 73 4092
rect -73 3832 -15 3844
rect -73 3526 -61 3832
rect -27 3526 -15 3832
rect -73 3514 -15 3526
rect 15 3832 73 3844
rect 15 3526 27 3832
rect 61 3526 73 3832
rect 15 3514 73 3526
rect -73 3266 -15 3278
rect -73 2960 -61 3266
rect -27 2960 -15 3266
rect -73 2948 -15 2960
rect 15 3266 73 3278
rect 15 2960 27 3266
rect 61 2960 73 3266
rect 15 2948 73 2960
rect -73 2700 -15 2712
rect -73 2394 -61 2700
rect -27 2394 -15 2700
rect -73 2382 -15 2394
rect 15 2700 73 2712
rect 15 2394 27 2700
rect 61 2394 73 2700
rect 15 2382 73 2394
rect -73 2134 -15 2146
rect -73 1828 -61 2134
rect -27 1828 -15 2134
rect -73 1816 -15 1828
rect 15 2134 73 2146
rect 15 1828 27 2134
rect 61 1828 73 2134
rect 15 1816 73 1828
rect -73 1568 -15 1580
rect -73 1262 -61 1568
rect -27 1262 -15 1568
rect -73 1250 -15 1262
rect 15 1568 73 1580
rect 15 1262 27 1568
rect 61 1262 73 1568
rect 15 1250 73 1262
rect -73 1002 -15 1014
rect -73 696 -61 1002
rect -27 696 -15 1002
rect -73 684 -15 696
rect 15 1002 73 1014
rect 15 696 27 1002
rect 61 696 73 1002
rect 15 684 73 696
rect -73 436 -15 448
rect -73 130 -61 436
rect -27 130 -15 436
rect -73 118 -15 130
rect 15 436 73 448
rect 15 130 27 436
rect 61 130 73 436
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -436 -61 -130
rect -27 -436 -15 -130
rect -73 -448 -15 -436
rect 15 -130 73 -118
rect 15 -436 27 -130
rect 61 -436 73 -130
rect 15 -448 73 -436
rect -73 -696 -15 -684
rect -73 -1002 -61 -696
rect -27 -1002 -15 -696
rect -73 -1014 -15 -1002
rect 15 -696 73 -684
rect 15 -1002 27 -696
rect 61 -1002 73 -696
rect 15 -1014 73 -1002
rect -73 -1262 -15 -1250
rect -73 -1568 -61 -1262
rect -27 -1568 -15 -1262
rect -73 -1580 -15 -1568
rect 15 -1262 73 -1250
rect 15 -1568 27 -1262
rect 61 -1568 73 -1262
rect 15 -1580 73 -1568
rect -73 -1828 -15 -1816
rect -73 -2134 -61 -1828
rect -27 -2134 -15 -1828
rect -73 -2146 -15 -2134
rect 15 -1828 73 -1816
rect 15 -2134 27 -1828
rect 61 -2134 73 -1828
rect 15 -2146 73 -2134
rect -73 -2394 -15 -2382
rect -73 -2700 -61 -2394
rect -27 -2700 -15 -2394
rect -73 -2712 -15 -2700
rect 15 -2394 73 -2382
rect 15 -2700 27 -2394
rect 61 -2700 73 -2394
rect 15 -2712 73 -2700
rect -73 -2960 -15 -2948
rect -73 -3266 -61 -2960
rect -27 -3266 -15 -2960
rect -73 -3278 -15 -3266
rect 15 -2960 73 -2948
rect 15 -3266 27 -2960
rect 61 -3266 73 -2960
rect 15 -3278 73 -3266
rect -73 -3526 -15 -3514
rect -73 -3832 -61 -3526
rect -27 -3832 -15 -3526
rect -73 -3844 -15 -3832
rect 15 -3526 73 -3514
rect 15 -3832 27 -3526
rect 61 -3832 73 -3526
rect 15 -3844 73 -3832
rect -73 -4092 -15 -4080
rect -73 -4398 -61 -4092
rect -27 -4398 -15 -4092
rect -73 -4410 -15 -4398
rect 15 -4092 73 -4080
rect 15 -4398 27 -4092
rect 61 -4398 73 -4092
rect 15 -4410 73 -4398
<< pdiffc >>
rect -61 4092 -27 4398
rect 27 4092 61 4398
rect -61 3526 -27 3832
rect 27 3526 61 3832
rect -61 2960 -27 3266
rect 27 2960 61 3266
rect -61 2394 -27 2700
rect 27 2394 61 2700
rect -61 1828 -27 2134
rect 27 1828 61 2134
rect -61 1262 -27 1568
rect 27 1262 61 1568
rect -61 696 -27 1002
rect 27 696 61 1002
rect -61 130 -27 436
rect 27 130 61 436
rect -61 -436 -27 -130
rect 27 -436 61 -130
rect -61 -1002 -27 -696
rect 27 -1002 61 -696
rect -61 -1568 -27 -1262
rect 27 -1568 61 -1262
rect -61 -2134 -27 -1828
rect 27 -2134 61 -1828
rect -61 -2700 -27 -2394
rect 27 -2700 61 -2394
rect -61 -3266 -27 -2960
rect 27 -3266 61 -2960
rect -61 -3832 -27 -3526
rect 27 -3832 61 -3526
rect -61 -4398 -27 -4092
rect 27 -4398 61 -4092
<< poly >>
rect -33 4491 33 4507
rect -33 4457 -17 4491
rect 17 4457 33 4491
rect -33 4441 33 4457
rect -15 4410 15 4441
rect -15 4049 15 4080
rect -33 4033 33 4049
rect -33 3999 -17 4033
rect 17 3999 33 4033
rect -33 3983 33 3999
rect -33 3925 33 3941
rect -33 3891 -17 3925
rect 17 3891 33 3925
rect -33 3875 33 3891
rect -15 3844 15 3875
rect -15 3483 15 3514
rect -33 3467 33 3483
rect -33 3433 -17 3467
rect 17 3433 33 3467
rect -33 3417 33 3433
rect -33 3359 33 3375
rect -33 3325 -17 3359
rect 17 3325 33 3359
rect -33 3309 33 3325
rect -15 3278 15 3309
rect -15 2917 15 2948
rect -33 2901 33 2917
rect -33 2867 -17 2901
rect 17 2867 33 2901
rect -33 2851 33 2867
rect -33 2793 33 2809
rect -33 2759 -17 2793
rect 17 2759 33 2793
rect -33 2743 33 2759
rect -15 2712 15 2743
rect -15 2351 15 2382
rect -33 2335 33 2351
rect -33 2301 -17 2335
rect 17 2301 33 2335
rect -33 2285 33 2301
rect -33 2227 33 2243
rect -33 2193 -17 2227
rect 17 2193 33 2227
rect -33 2177 33 2193
rect -15 2146 15 2177
rect -15 1785 15 1816
rect -33 1769 33 1785
rect -33 1735 -17 1769
rect 17 1735 33 1769
rect -33 1719 33 1735
rect -33 1661 33 1677
rect -33 1627 -17 1661
rect 17 1627 33 1661
rect -33 1611 33 1627
rect -15 1580 15 1611
rect -15 1219 15 1250
rect -33 1203 33 1219
rect -33 1169 -17 1203
rect 17 1169 33 1203
rect -33 1153 33 1169
rect -33 1095 33 1111
rect -33 1061 -17 1095
rect 17 1061 33 1095
rect -33 1045 33 1061
rect -15 1014 15 1045
rect -15 653 15 684
rect -33 637 33 653
rect -33 603 -17 637
rect 17 603 33 637
rect -33 587 33 603
rect -33 529 33 545
rect -33 495 -17 529
rect 17 495 33 529
rect -33 479 33 495
rect -15 448 15 479
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -479 15 -448
rect -33 -495 33 -479
rect -33 -529 -17 -495
rect 17 -529 33 -495
rect -33 -545 33 -529
rect -33 -603 33 -587
rect -33 -637 -17 -603
rect 17 -637 33 -603
rect -33 -653 33 -637
rect -15 -684 15 -653
rect -15 -1045 15 -1014
rect -33 -1061 33 -1045
rect -33 -1095 -17 -1061
rect 17 -1095 33 -1061
rect -33 -1111 33 -1095
rect -33 -1169 33 -1153
rect -33 -1203 -17 -1169
rect 17 -1203 33 -1169
rect -33 -1219 33 -1203
rect -15 -1250 15 -1219
rect -15 -1611 15 -1580
rect -33 -1627 33 -1611
rect -33 -1661 -17 -1627
rect 17 -1661 33 -1627
rect -33 -1677 33 -1661
rect -33 -1735 33 -1719
rect -33 -1769 -17 -1735
rect 17 -1769 33 -1735
rect -33 -1785 33 -1769
rect -15 -1816 15 -1785
rect -15 -2177 15 -2146
rect -33 -2193 33 -2177
rect -33 -2227 -17 -2193
rect 17 -2227 33 -2193
rect -33 -2243 33 -2227
rect -33 -2301 33 -2285
rect -33 -2335 -17 -2301
rect 17 -2335 33 -2301
rect -33 -2351 33 -2335
rect -15 -2382 15 -2351
rect -15 -2743 15 -2712
rect -33 -2759 33 -2743
rect -33 -2793 -17 -2759
rect 17 -2793 33 -2759
rect -33 -2809 33 -2793
rect -33 -2867 33 -2851
rect -33 -2901 -17 -2867
rect 17 -2901 33 -2867
rect -33 -2917 33 -2901
rect -15 -2948 15 -2917
rect -15 -3309 15 -3278
rect -33 -3325 33 -3309
rect -33 -3359 -17 -3325
rect 17 -3359 33 -3325
rect -33 -3375 33 -3359
rect -33 -3433 33 -3417
rect -33 -3467 -17 -3433
rect 17 -3467 33 -3433
rect -33 -3483 33 -3467
rect -15 -3514 15 -3483
rect -15 -3875 15 -3844
rect -33 -3891 33 -3875
rect -33 -3925 -17 -3891
rect 17 -3925 33 -3891
rect -33 -3941 33 -3925
rect -33 -3999 33 -3983
rect -33 -4033 -17 -3999
rect 17 -4033 33 -3999
rect -33 -4049 33 -4033
rect -15 -4080 15 -4049
rect -15 -4441 15 -4410
rect -33 -4457 33 -4441
rect -33 -4491 -17 -4457
rect 17 -4491 33 -4457
rect -33 -4507 33 -4491
<< polycont >>
rect -17 4457 17 4491
rect -17 3999 17 4033
rect -17 3891 17 3925
rect -17 3433 17 3467
rect -17 3325 17 3359
rect -17 2867 17 2901
rect -17 2759 17 2793
rect -17 2301 17 2335
rect -17 2193 17 2227
rect -17 1735 17 1769
rect -17 1627 17 1661
rect -17 1169 17 1203
rect -17 1061 17 1095
rect -17 603 17 637
rect -17 495 17 529
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -529 17 -495
rect -17 -637 17 -603
rect -17 -1095 17 -1061
rect -17 -1203 17 -1169
rect -17 -1661 17 -1627
rect -17 -1769 17 -1735
rect -17 -2227 17 -2193
rect -17 -2335 17 -2301
rect -17 -2793 17 -2759
rect -17 -2901 17 -2867
rect -17 -3359 17 -3325
rect -17 -3467 17 -3433
rect -17 -3925 17 -3891
rect -17 -4033 17 -3999
rect -17 -4491 17 -4457
<< locali >>
rect -33 4457 -17 4491
rect 17 4457 33 4491
rect -61 4398 -27 4414
rect -61 4076 -27 4092
rect 27 4398 61 4414
rect 27 4076 61 4092
rect -33 3999 -17 4033
rect 17 3999 33 4033
rect -33 3891 -17 3925
rect 17 3891 33 3925
rect -61 3832 -27 3848
rect -61 3510 -27 3526
rect 27 3832 61 3848
rect 27 3510 61 3526
rect -33 3433 -17 3467
rect 17 3433 33 3467
rect -33 3325 -17 3359
rect 17 3325 33 3359
rect -61 3266 -27 3282
rect -61 2944 -27 2960
rect 27 3266 61 3282
rect 27 2944 61 2960
rect -33 2867 -17 2901
rect 17 2867 33 2901
rect -33 2759 -17 2793
rect 17 2759 33 2793
rect -61 2700 -27 2716
rect -61 2378 -27 2394
rect 27 2700 61 2716
rect 27 2378 61 2394
rect -33 2301 -17 2335
rect 17 2301 33 2335
rect -33 2193 -17 2227
rect 17 2193 33 2227
rect -61 2134 -27 2150
rect -61 1812 -27 1828
rect 27 2134 61 2150
rect 27 1812 61 1828
rect -33 1735 -17 1769
rect 17 1735 33 1769
rect -33 1627 -17 1661
rect 17 1627 33 1661
rect -61 1568 -27 1584
rect -61 1246 -27 1262
rect 27 1568 61 1584
rect 27 1246 61 1262
rect -33 1169 -17 1203
rect 17 1169 33 1203
rect -33 1061 -17 1095
rect 17 1061 33 1095
rect -61 1002 -27 1018
rect -61 680 -27 696
rect 27 1002 61 1018
rect 27 680 61 696
rect -33 603 -17 637
rect 17 603 33 637
rect -33 495 -17 529
rect 17 495 33 529
rect -61 436 -27 452
rect -61 114 -27 130
rect 27 436 61 452
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -452 -27 -436
rect 27 -130 61 -114
rect 27 -452 61 -436
rect -33 -529 -17 -495
rect 17 -529 33 -495
rect -33 -637 -17 -603
rect 17 -637 33 -603
rect -61 -696 -27 -680
rect -61 -1018 -27 -1002
rect 27 -696 61 -680
rect 27 -1018 61 -1002
rect -33 -1095 -17 -1061
rect 17 -1095 33 -1061
rect -33 -1203 -17 -1169
rect 17 -1203 33 -1169
rect -61 -1262 -27 -1246
rect -61 -1584 -27 -1568
rect 27 -1262 61 -1246
rect 27 -1584 61 -1568
rect -33 -1661 -17 -1627
rect 17 -1661 33 -1627
rect -33 -1769 -17 -1735
rect 17 -1769 33 -1735
rect -61 -1828 -27 -1812
rect -61 -2150 -27 -2134
rect 27 -1828 61 -1812
rect 27 -2150 61 -2134
rect -33 -2227 -17 -2193
rect 17 -2227 33 -2193
rect -33 -2335 -17 -2301
rect 17 -2335 33 -2301
rect -61 -2394 -27 -2378
rect -61 -2716 -27 -2700
rect 27 -2394 61 -2378
rect 27 -2716 61 -2700
rect -33 -2793 -17 -2759
rect 17 -2793 33 -2759
rect -33 -2901 -17 -2867
rect 17 -2901 33 -2867
rect -61 -2960 -27 -2944
rect -61 -3282 -27 -3266
rect 27 -2960 61 -2944
rect 27 -3282 61 -3266
rect -33 -3359 -17 -3325
rect 17 -3359 33 -3325
rect -33 -3467 -17 -3433
rect 17 -3467 33 -3433
rect -61 -3526 -27 -3510
rect -61 -3848 -27 -3832
rect 27 -3526 61 -3510
rect 27 -3848 61 -3832
rect -33 -3925 -17 -3891
rect 17 -3925 33 -3891
rect -33 -4033 -17 -3999
rect 17 -4033 33 -3999
rect -61 -4092 -27 -4076
rect -61 -4414 -27 -4398
rect 27 -4092 61 -4076
rect 27 -4414 61 -4398
rect -33 -4491 -17 -4457
rect 17 -4491 33 -4457
<< viali >>
rect -17 4457 17 4491
rect -61 4092 -27 4398
rect 27 4092 61 4398
rect -17 3999 17 4033
rect -17 3891 17 3925
rect -61 3526 -27 3832
rect 27 3526 61 3832
rect -17 3433 17 3467
rect -17 3325 17 3359
rect -61 2960 -27 3266
rect 27 2960 61 3266
rect -17 2867 17 2901
rect -17 2759 17 2793
rect -61 2394 -27 2700
rect 27 2394 61 2700
rect -17 2301 17 2335
rect -17 2193 17 2227
rect -61 1828 -27 2134
rect 27 1828 61 2134
rect -17 1735 17 1769
rect -17 1627 17 1661
rect -61 1262 -27 1568
rect 27 1262 61 1568
rect -17 1169 17 1203
rect -17 1061 17 1095
rect -61 696 -27 1002
rect 27 696 61 1002
rect -17 603 17 637
rect -17 495 17 529
rect -61 130 -27 436
rect 27 130 61 436
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -436 -27 -130
rect 27 -436 61 -130
rect -17 -529 17 -495
rect -17 -637 17 -603
rect -61 -1002 -27 -696
rect 27 -1002 61 -696
rect -17 -1095 17 -1061
rect -17 -1203 17 -1169
rect -61 -1568 -27 -1262
rect 27 -1568 61 -1262
rect -17 -1661 17 -1627
rect -17 -1769 17 -1735
rect -61 -2134 -27 -1828
rect 27 -2134 61 -1828
rect -17 -2227 17 -2193
rect -17 -2335 17 -2301
rect -61 -2700 -27 -2394
rect 27 -2700 61 -2394
rect -17 -2793 17 -2759
rect -17 -2901 17 -2867
rect -61 -3266 -27 -2960
rect 27 -3266 61 -2960
rect -17 -3359 17 -3325
rect -17 -3467 17 -3433
rect -61 -3832 -27 -3526
rect 27 -3832 61 -3526
rect -17 -3925 17 -3891
rect -17 -4033 17 -3999
rect -61 -4398 -27 -4092
rect 27 -4398 61 -4092
rect -17 -4491 17 -4457
<< metal1 >>
rect -29 4491 29 4497
rect -29 4457 -17 4491
rect 17 4457 29 4491
rect -29 4451 29 4457
rect -67 4398 -21 4410
rect -67 4092 -61 4398
rect -27 4092 -21 4398
rect -67 4080 -21 4092
rect 21 4398 67 4410
rect 21 4092 27 4398
rect 61 4092 67 4398
rect 21 4080 67 4092
rect -29 4033 29 4039
rect -29 3999 -17 4033
rect 17 3999 29 4033
rect -29 3993 29 3999
rect -29 3925 29 3931
rect -29 3891 -17 3925
rect 17 3891 29 3925
rect -29 3885 29 3891
rect -67 3832 -21 3844
rect -67 3526 -61 3832
rect -27 3526 -21 3832
rect -67 3514 -21 3526
rect 21 3832 67 3844
rect 21 3526 27 3832
rect 61 3526 67 3832
rect 21 3514 67 3526
rect -29 3467 29 3473
rect -29 3433 -17 3467
rect 17 3433 29 3467
rect -29 3427 29 3433
rect -29 3359 29 3365
rect -29 3325 -17 3359
rect 17 3325 29 3359
rect -29 3319 29 3325
rect -67 3266 -21 3278
rect -67 2960 -61 3266
rect -27 2960 -21 3266
rect -67 2948 -21 2960
rect 21 3266 67 3278
rect 21 2960 27 3266
rect 61 2960 67 3266
rect 21 2948 67 2960
rect -29 2901 29 2907
rect -29 2867 -17 2901
rect 17 2867 29 2901
rect -29 2861 29 2867
rect -29 2793 29 2799
rect -29 2759 -17 2793
rect 17 2759 29 2793
rect -29 2753 29 2759
rect -67 2700 -21 2712
rect -67 2394 -61 2700
rect -27 2394 -21 2700
rect -67 2382 -21 2394
rect 21 2700 67 2712
rect 21 2394 27 2700
rect 61 2394 67 2700
rect 21 2382 67 2394
rect -29 2335 29 2341
rect -29 2301 -17 2335
rect 17 2301 29 2335
rect -29 2295 29 2301
rect -29 2227 29 2233
rect -29 2193 -17 2227
rect 17 2193 29 2227
rect -29 2187 29 2193
rect -67 2134 -21 2146
rect -67 1828 -61 2134
rect -27 1828 -21 2134
rect -67 1816 -21 1828
rect 21 2134 67 2146
rect 21 1828 27 2134
rect 61 1828 67 2134
rect 21 1816 67 1828
rect -29 1769 29 1775
rect -29 1735 -17 1769
rect 17 1735 29 1769
rect -29 1729 29 1735
rect -29 1661 29 1667
rect -29 1627 -17 1661
rect 17 1627 29 1661
rect -29 1621 29 1627
rect -67 1568 -21 1580
rect -67 1262 -61 1568
rect -27 1262 -21 1568
rect -67 1250 -21 1262
rect 21 1568 67 1580
rect 21 1262 27 1568
rect 61 1262 67 1568
rect 21 1250 67 1262
rect -29 1203 29 1209
rect -29 1169 -17 1203
rect 17 1169 29 1203
rect -29 1163 29 1169
rect -29 1095 29 1101
rect -29 1061 -17 1095
rect 17 1061 29 1095
rect -29 1055 29 1061
rect -67 1002 -21 1014
rect -67 696 -61 1002
rect -27 696 -21 1002
rect -67 684 -21 696
rect 21 1002 67 1014
rect 21 696 27 1002
rect 61 696 67 1002
rect 21 684 67 696
rect -29 637 29 643
rect -29 603 -17 637
rect 17 603 29 637
rect -29 597 29 603
rect -29 529 29 535
rect -29 495 -17 529
rect 17 495 29 529
rect -29 489 29 495
rect -67 436 -21 448
rect -67 130 -61 436
rect -27 130 -21 436
rect -67 118 -21 130
rect 21 436 67 448
rect 21 130 27 436
rect 61 130 67 436
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -436 -61 -130
rect -27 -436 -21 -130
rect -67 -448 -21 -436
rect 21 -130 67 -118
rect 21 -436 27 -130
rect 61 -436 67 -130
rect 21 -448 67 -436
rect -29 -495 29 -489
rect -29 -529 -17 -495
rect 17 -529 29 -495
rect -29 -535 29 -529
rect -29 -603 29 -597
rect -29 -637 -17 -603
rect 17 -637 29 -603
rect -29 -643 29 -637
rect -67 -696 -21 -684
rect -67 -1002 -61 -696
rect -27 -1002 -21 -696
rect -67 -1014 -21 -1002
rect 21 -696 67 -684
rect 21 -1002 27 -696
rect 61 -1002 67 -696
rect 21 -1014 67 -1002
rect -29 -1061 29 -1055
rect -29 -1095 -17 -1061
rect 17 -1095 29 -1061
rect -29 -1101 29 -1095
rect -29 -1169 29 -1163
rect -29 -1203 -17 -1169
rect 17 -1203 29 -1169
rect -29 -1209 29 -1203
rect -67 -1262 -21 -1250
rect -67 -1568 -61 -1262
rect -27 -1568 -21 -1262
rect -67 -1580 -21 -1568
rect 21 -1262 67 -1250
rect 21 -1568 27 -1262
rect 61 -1568 67 -1262
rect 21 -1580 67 -1568
rect -29 -1627 29 -1621
rect -29 -1661 -17 -1627
rect 17 -1661 29 -1627
rect -29 -1667 29 -1661
rect -29 -1735 29 -1729
rect -29 -1769 -17 -1735
rect 17 -1769 29 -1735
rect -29 -1775 29 -1769
rect -67 -1828 -21 -1816
rect -67 -2134 -61 -1828
rect -27 -2134 -21 -1828
rect -67 -2146 -21 -2134
rect 21 -1828 67 -1816
rect 21 -2134 27 -1828
rect 61 -2134 67 -1828
rect 21 -2146 67 -2134
rect -29 -2193 29 -2187
rect -29 -2227 -17 -2193
rect 17 -2227 29 -2193
rect -29 -2233 29 -2227
rect -29 -2301 29 -2295
rect -29 -2335 -17 -2301
rect 17 -2335 29 -2301
rect -29 -2341 29 -2335
rect -67 -2394 -21 -2382
rect -67 -2700 -61 -2394
rect -27 -2700 -21 -2394
rect -67 -2712 -21 -2700
rect 21 -2394 67 -2382
rect 21 -2700 27 -2394
rect 61 -2700 67 -2394
rect 21 -2712 67 -2700
rect -29 -2759 29 -2753
rect -29 -2793 -17 -2759
rect 17 -2793 29 -2759
rect -29 -2799 29 -2793
rect -29 -2867 29 -2861
rect -29 -2901 -17 -2867
rect 17 -2901 29 -2867
rect -29 -2907 29 -2901
rect -67 -2960 -21 -2948
rect -67 -3266 -61 -2960
rect -27 -3266 -21 -2960
rect -67 -3278 -21 -3266
rect 21 -2960 67 -2948
rect 21 -3266 27 -2960
rect 61 -3266 67 -2960
rect 21 -3278 67 -3266
rect -29 -3325 29 -3319
rect -29 -3359 -17 -3325
rect 17 -3359 29 -3325
rect -29 -3365 29 -3359
rect -29 -3433 29 -3427
rect -29 -3467 -17 -3433
rect 17 -3467 29 -3433
rect -29 -3473 29 -3467
rect -67 -3526 -21 -3514
rect -67 -3832 -61 -3526
rect -27 -3832 -21 -3526
rect -67 -3844 -21 -3832
rect 21 -3526 67 -3514
rect 21 -3832 27 -3526
rect 61 -3832 67 -3526
rect 21 -3844 67 -3832
rect -29 -3891 29 -3885
rect -29 -3925 -17 -3891
rect 17 -3925 29 -3891
rect -29 -3931 29 -3925
rect -29 -3999 29 -3993
rect -29 -4033 -17 -3999
rect 17 -4033 29 -3999
rect -29 -4039 29 -4033
rect -67 -4092 -21 -4080
rect -67 -4398 -61 -4092
rect -27 -4398 -21 -4092
rect -67 -4410 -21 -4398
rect 21 -4092 67 -4080
rect 21 -4398 27 -4092
rect 61 -4398 67 -4092
rect 21 -4410 67 -4398
rect -29 -4457 29 -4451
rect -29 -4491 -17 -4457
rect 17 -4491 29 -4457
rect -29 -4497 29 -4491
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.65 l 0.15 m 16 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
