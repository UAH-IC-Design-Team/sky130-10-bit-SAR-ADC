magic
tech sky130A
magscale 1 2
timestamp 1668103091
<< error_s >>
rect -5706188 -6573006 -5706160 -6572950
rect -5706132 -6573006 -5706104 -6572950
rect -5706515 -6577297 -5706315 -6577245
rect -5706195 -6577297 -5706065 -6577245
rect -5706515 -6577381 -5706315 -6577327
rect -5706195 -6577381 -5706065 -6577327
rect -5706515 -6577463 -5706315 -6577411
rect -5706195 -6577463 -5706065 -6577411
<< metal1 >>
rect -5841100 -6572040 -5837740 -6572020
rect -5841100 -6572420 -5838140 -6572040
rect -5837760 -6572420 -5837740 -6572040
rect -5841100 -6572440 -5837740 -6572420
rect -5841100 -6572820 -5837740 -6572800
rect -5841100 -6573200 -5838140 -6572820
rect -5837760 -6573200 -5837740 -6572820
rect -5841100 -6573220 -5837740 -6573200
<< via1 >>
rect -5838140 -6572420 -5837760 -6572040
rect -5838140 -6573200 -5837760 -6572820
<< metal2 >>
rect -5838160 -6571120 -5837740 -6571100
rect -5838160 -6571480 -5838140 -6571120
rect -5837760 -6571480 -5837740 -6571120
rect -5838160 -6572040 -5837740 -6571480
rect -5838160 -6572420 -5838140 -6572040
rect -5837760 -6572420 -5837740 -6572040
rect -5838160 -6572440 -5837740 -6572420
rect -5838160 -6572820 -5837740 -6572800
rect -5838160 -6573200 -5838140 -6572820
rect -5837760 -6573200 -5837740 -6572820
rect -5838160 -6573720 -5837740 -6573200
rect -5838160 -6574080 -5838140 -6573720
rect -5837760 -6574080 -5837740 -6573720
rect -5838160 -6574100 -5837740 -6574080
<< via2 >>
rect -5838140 -6571480 -5837760 -6571120
rect -5838140 -6574080 -5837760 -6573720
<< metal3 >>
rect -5838160 -6571120 -5837740 -6571100
rect -5838160 -6571480 -5838140 -6571120
rect -5837760 -6571480 -5837740 -6571120
rect -5838160 -6571500 -5837740 -6571480
rect -5838160 -6573720 -5837740 -6573700
rect -5838160 -6574080 -5838140 -6573720
rect -5837760 -6574080 -5837740 -6573720
rect -5838160 -6574100 -5837740 -6574080
<< via3 >>
rect -5838140 -6571480 -5837760 -6571120
rect -5838140 -6574080 -5837760 -6573720
<< metal4 >>
rect -5838160 -6571120 -5716380 -6571100
rect -5838160 -6571480 -5838140 -6571120
rect -5837760 -6571480 -5716380 -6571120
rect -5838160 -6571500 -5716380 -6571480
rect -5838160 -6573720 -5716380 -6573700
rect -5838160 -6574080 -5838140 -6573720
rect -5837760 -6574080 -5716380 -6573720
rect -5838160 -6574100 -5716380 -6574080
use bootstrapped_sampling_switch  bootstrapped_sampling_switch_0
timestamp 1667491297
transform 0 1 -5836200 -1 0 -6565850
box -3600 -5100 17150 2800
use comparator  comparator_0
timestamp 1668055187
transform 0 -1 -5701200 1 0 -6584490
box 6930 4070 16410 8800
use controller  controller_0 OpenLane/designs/controller/runs/RUN_2022.11.08_16.38.24/results/final/mag
timestamp 1668055187
transform 1 0 -5704000 0 1 -6585000
box 0 0 21861 24005
use dac  dac_0
timestamp 1668103091
transform 1 0 -5798000 0 1 -6624400
box -35000 33000 88200 70300
<< end >>
